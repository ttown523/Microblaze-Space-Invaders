XlxV64EB    5cd2    1440�ݥ��.�Rʅ�T^�b�5a�o�hL4��O��������ν�"�o�p!�'�q�._U�F�$��85�3o=��n�]0�}��&y��ƾ������
�Fxe{��AwvY��w
~	�_Ӯ8���N@:�;��r�?ktV�"��L�k^Y(A�����\Im��$4u�h�R���4ҨG��G���N��S�����ķ�`J�uQ_��U>�j��Z��]���8�n�*�W�֐@���W��507N�#;f�+�*�^<u
|�_-�ě�WT�E�G��r5��	�h�d��X;a�rѲ���D���Y�!���Q9��;o��A��}y��k�a�Ԣ0��j��W���NC�gEi���4�TE��q����dh�K�ۋ�ϐj�h\��c��u�sQ�(��`t�_-��T��T2f�������0�m]F{؊)M�W�^5���!�>XT�p�J0া�	�6f;�ߢm����S0%x:2��F,��4���[������7�g�/���ne�s��_��+�ֵG�����9�b-�R��7�z�nJ�4�H�;&�\�8L�G~e�ʕl�W��{a"�[��J�ʆ��+�������_PSń��C���>;x16,A�|\M3wM�~��̥��@"~U�>��Y]/Qta{χ����5�B��ش�oO/��6��l��Y^% jQ%����s���n���vJ�I�c�:/������?�l�9����i�I���E�fe]Z�B?t)=��%�J����d��_��]�Q�<�1ȥ�k;1-�Ri��1f��Sm|k.��l�{^���C�h#xw�q��4����M��J2K��s<c��v�t�n�j�<�\��n��:�VK���\krv~��o-K�^H��]�c�M�^
Gy
|�~Z�5g����#�1�t����Җ�4d��9Gb�L�/_@�!�m��&�j�HQgF��I�Ϲ[�7�*��v��k�SPR}����9A�N`�@Ɓ��0��k:U�+
큰~�[���\�,p�~�HS6�f��S����p$��"������Y�H�..|�Y�`��fɴ(�����@6�ɐ���'�I��H>x{M 5��Cfzv{��j��^!�x��Z��70u_"WlR%������z~�ԫ4�39e�9�v¡��Qp�@���S��j�t�e$�8��Tż���O�4��j}���	�੭���
���~F�cQ�Ts���0r����O�����]/���&�{���%��n�^_���*�tVy�n٧��We��x8ް�a9�ķ���-dL<��I���~E����~:$�eήق#m���\�CK���]PD�Y�	�&�ܔ��j�a�JU��c�C�	+�w#��?�Q�oB*�� {�f�[�P��ᵍOp�`5���W�v{7��wb��D˲��Z��r
c�a���0,���	�P��x�{��"ļ�@yE'D��B�8@��ߞ�y'CхNH�����3ϷBV/�Y��]�3A�v�]�ʣ�����X%l*Ԃ�=0�&���˒6H��R������q{��BߚT��4l��r<�}*d��i��"�:k]�w��z^�Ӓ\o�u��r�3`�#��%�h[����Fښ9t�Udރ���#N���F?a0��%�
�����T&.K/��>���l�t+y"�)%.�F!")է���}Dɝ?�s�����
J�5�b����d�C~��s�y�J����������SiO]�ߴ�cbJ��kC�S��aɅ{p[��dX�����{��H��d��G�� : ����0"uQ�8q1{lc��ۥy��Ĩ���l�:٭���Rc]�D	lN���*{��c����(
0ǽ�����J�Ev,��'U,!��h�$��Q�N��{{P<f�Fם!͟@%sq*'��q�5�d�V�`�x1���Ȱ��K]�@������G�����A�%W��Й�/���PV����Dȇaؤ��H��s���@v��%>p��nP��-a�Z�N�m�T��vj�U�X8p��3���؍']1�Xקo(յ���G`�'�� !)O�t7`/�ٶ;ï:�c(���i��Z��&5�#H����|��,I\�N��O[y����\z@�h9�ށi�M�Ӧߌ�����}j�*���cC��%k,#L���ʀ��!h������omW�utRNkJ�(ղ��a���6)�����xhԍ�[���e�;n(�%�D�H����8;�>T곇+���^}]������gT��v|y7�z�����W��A�̃Vzed�r���>���ix�J9�Z�������L�k�h\a�Āe3wK�VS��<�R6���<�]o����lB۬v��i�$��(�-t�s�=M!������LJ�
�����c�I��(����i�F�tѡ?2pQ=�LxZX��l����߼y�K�
�����H�r+�|a:�S��İ��#�~'K_��B�w�)�)�����ج��j�8U��^�� �Ƶ}�x�;�
H����>�/u���'�G[ B��gK�̗�M��]��%N�Q�.���՛��~���MNև�p�P�x����)(��C���EBxXaNv8ݨҙ�a��z��V^�U
Kߛ�����)#�u����Ǐd'Ekg��=�Zb��;_�!Ha4��*1Y=۠ӊ��:|�L�-�C%��V��q�}���T��8��*#�右:a'�5
���x}�܄ͬ�F
�z�q�R4$���p-��i^�A�U���(վ�B�b����B>�n j�2��I�
x\8���D�x�]`��ݹ�xY�6&��B�R��9�)h(}������p�#SѢ�8Wrf3:l�d4�I�q�x�q�gv�P�KU����란Yt��㻙\�++ѱ�I��5�����k�[�k-$�����!�B�<�'���ܺ�c�F#7�#f?�d�������H!��)!R	������ ��N�z�m!��br����K��m;9$"2����XSZ��:�D�\�1�#o��o�*	�ͳ^Ԣ�q�#ˠ��a}�ƏJ]��Dw�M�\rm�v�Y�d<�*-u�<r�͎���L�����|Roϑ}7bt{�Ө�P#����lf���˲7Ľ���S�ﳨ�͗��n��fK���F�?�ꄵT����$�s�vZ:�2m�cm(����廮�c��_���[�I��tO�d���%/��9_'�?��4��r_��,�/Z�&�x�G@�j�R���'�㬌_p�S�qR��7�TCҀ�̯)�Лz�'�mK���Q�G����;��ZiK7���E����T)M3ΓNY�~�lI5=��C����f���]�/yJ�b�%��.��D�wv3Fx^���go��ӓzT��>8�8��h�ܱ���<�4�����h�B�ъ.r_���ux�V n� �i矟��������1���˶��[�.���o���Ʊ���\'����}k�\�%���*��B�S��bj�$<ą0���o��̱h ��!��C�Ovk����
K��pޯ�
����pCa�� �P��	�[�:1�or�2�S�,�ᙾLA(�9���8�[$��8�ڋ�z"�G�P������@�o��o�{� S|5z��cQ]�o����u�>� F�.xޖ�� ������YC��/@_���%��G�畚o@�D!e�s���L�>qz?i�i{a_���/,ZBu�X���e1�2Dc�<��6� i�D��.�h��S�C��:���;�J���_��o�{݁R�����u�\������o��G�-^6n�����k��kF��S�2V��pT��u�tfT�sJJwx75�U8v�G�N���ᒾz�e�P{شi0)��'���1�|ɞG�d�����P
\��%�J�1 ��v3�!��'nȾc���*yg�����yԯEi�����/'q!QIr� ����_�۔א��;6�l��7���.R�@i����M���>$BZy� ��q4<@���R�.-��9T�U� ��H5����c�׸Ǵ�*�\�#%�O� Wd����=D]�bw!���J �0+��!��R��wӠ��8�Ȁ?c0����M�/1�+C&P�y'	� z+K����x���4��[K�K��00P��-��_���F�S�l�i}:gZG�����L��k:��w��gOq����g���A�3ς|r��I(�\Op��z��K
.�:�C}*��7������i��AFiۛM�t����>@M����'�4�`�h�H���3طcC��I����E|�m6o%O�n-n��1���n�l�%��aɝ֬�Ԗ�\�c��y��lR�����Qy^����3]T�ȐT�\�#\(��ή��$�8� >5�$Y�����oz8��d�g-E���d���H�H�{V��wsd��~�).gQ��kݳ��
��sY��6�^p�d=s�������	�4�@�5�����*+0[
;����S+-��Ψ��"n\>�0���f`��Ϻx8Z$����%ٞ�����`g�|��=e�6Ĉ-f��R�O����[���Y���rIik�$�dA,����$�G�5*�4[��Ų�Uj%����^�/Mf� ǣ�������1�`�"i��XRJ0���U]f�`z0,N�����������D��q$��b�������D�=���� `(Wi����������W(A�sE9�Tј�J��ț�I/����|D�/��jzK��KG�=c������-���}:N:]���WZ�%���g��3WWp������
��6�;+oZ>�]�u=P�@�7�^屝�����(#� (	�f�@�
���/��Y��^�g����!m��lT��Y1���jK'�5�O�D��r�Z����?��"���N,u������S"�zq���TNv,��	� ~��Ɣ#�!F�{�,%���=�@���	�U���,!2�twf?'H�H�⤽��e��m#b�Y�_��
9�԰|��O��? �� �Źtdia:<W෪��$
��ʐ�9y.g���������H������ٜ�^�8