XlxV64EB    2e8b     cc0��:�܌�G���o��nf@@��Y��.7Y#�_S��9��!���+3��h�n^}�D��J`��T$}9.ȠV`�*F$�b�7S{��3�nXzڿ<�^�������T�i�B������{�5��3�ߵ.�)c��� s+0ʹ�8a,	���/���JR�a/ ��'�f��~��3�-��K�
��ep���}f�I���^H�8\��M(��%9�a:��Fʼ��!��)��1♊k��6H�/���_>t�B۩�'#�L�|�8��j��2��Ŀ`����N<ʼ.��M����B�@�ḵ��x��K��(G4�?�N}v6�eΕ�\�&��S]dҕ��ŐFw�$Ғw�"<��1���FaMk�wn���#��&���S��T'%�����ݕ��|�^������u�6!Z�!��9�uz��U<�����UL��b��dGMa@���♋oЌ
Ӣ���Eh;��/��{ar�!�u*)����A��R�]F��c�ߐ�]�5�Ȝ�|%_+���#jY�6܇�E��~2k,0��X�,<����ʌ3rGWQ���Ӆk�.�:�@�.J�?�1BCKI�����e"*��S�nR{9bk�cf�� 5��KAi�����D)oj�� �,ԷK��9��e�Kd����n`�)9Q����u8ӵe��Q�UHˁԋ}u��'���Ĩ�߂ �_P_s��k�nP3�4U��u��r��{�7��i(����b�(3�k�^O�QSş�Q��~d���r���W_�GK5/Tҳ�OnS�̯�"{r$��7��b��tGa�b5�6` -�fq��}��K�n}��>�������5Ȓ����3k]y�g�ڈ  ��֭q��y��D��^�n_~��c;ƬK0�S�mV���,�x��n}����F����Gv����٣m������9&x���߯T2�/��Lim������/��Jt]S��AM��\|���ԯ%d����m-�� bEaZ�zw��*� 5(Z��bZ��S2ka�9k:V0��u��3gǯ"~H߲4�b^".k��9�t�F�F�!O��r���KB�T=ן3|���#-����X.��Z�[+9WTf��6� �0�]  ���2�i��"�Hl�\ɇӷ���ߴ?"��',V@i�G�7*|�`gO��(c����UB�	6��^y��:e? _��@$q�ӥ�R��t��|lz+���	ǅ_դ�J��a	���QC��� r'��ِ^L6c����9���_]����%n�y \�{z䐪@P�!lף+�E�ˈ���s��Z����`�)���W߀��ǧ�8���Z7����O�B,Z��]w]@O��H&�������x$��U{���e�\��Б,<�ި'�A7�0e�V������t6�@z&��I�̮LIaП��!R���D���\r�5s`J;�c�3̺����9\��؛=�&#Z�6��5JV���>Le�<=}=S��я6�ړ���EaUm� #P�	s���o�`�>�_	�ԑ����vi��>��Z%��C�K?ۘ�,9���S��z��q���<��P�&J>у���R��&e�䪝�zYNC<g�B1��+�(�T:�e��~��!@�h�<����CЙklb�J�}���$}��������/cHE2����~�r�V���9��]z\�Wn��7=&�Z?�dՋ'����V��r��W�����[�?�%o�2��K�l�"N��]YKv:�Ҧ(vO
������px	]EE�-�Q^�>��R>���`�YS�W��.�j�,4]-&N:�<�x��=~��ei7<l3�f�3j�eأ��RH��c�R��c{��p�5+<���"���`�����F�hA�{��������N��2dy��
!w%��8����(ѶB�d�3"��b����u6|%j|�"�wU3A����b�k��QÓ�w]���H(�T���S�y��$8}�8�
|�W��. ��NQc/HV�U���֔;D�!�-Fq>+��3���PH��Э��enq�$w�B"Nw��ÛY��)���\��������L����s�3N{;�k]BF鉀������3��@�mu�^��d��]nj��ﻏ�F���}/N�Śe�p=Rx�d�2JhyL�|G�7@��h`c�R�=��ot$�����X� �,E��s/bxQ��n��Rd%c��J��G*S�5T�3��c�6�j�9Q0�goyϾ��t8�E�U��71g�V*�!���c�����&�[��� �T��%���tu6��� F��%���e_k���	��9 �j�`I3��?���j�o����������%7�Gx��88� `V&��ʿw͗����I�#wB��@y�Ӵ��Uƍ�4R~���&�7Y���p�
������WrF���BS֍ګ���������N�j��G�nE�T���;��OSef��R|��8`����go���E]w�����:��l�I�惻�>̼��X�al�~�@�}��p$pZ*��H*lu`IX���_=t{W�܉Y����C��`�>?���r�;�;5[���p�ݐ%M".=}fV�VѴ5m*f��O�]��K�K�&���nC�C���`�V�ʽ~q��ކ0Zeںj��L��Eg|hN�s!�6e��iń)`�2E�a�����H���;�ǋ�:g�<�P�Y���-��<�[���/�P�KZz�Rk�+�$&���1G_��,���[m
0��x������)�����p	6;�ë��3��<�t'dc�3�������� DjF�/v���v����p�}���GTl.9&�&~�Í�Č�u���pmؖw�Y���%Σ��5N��ˢ�4�;���3ݞ���8�g��Cl�	�!��=SOKR���RBTw1� ��b��Z�Ii�A�fw�xiU�sog��3
iPEF�H*���M,4�[Pix�`�$�sr�D��_������ZNr�u��<#zS��S�����&g+v���ʭ͚�s��s�'P��~��?K"^��NY��E�I"�ڭ�C�1ك\��ÀݕlL� W65�o~���E&�r}�`gq��"bj`����ۘ��Թ� 9q#V	WGJ��n}����"1u�� -��Nvѡ���}U2�#��]zqF���CiK!K�����A�&E&$aO_�g�	��t_J$7#i�����a ���e�