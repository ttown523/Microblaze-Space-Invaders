XlxV64EB    fa00    2d10c���c�+FD&�Ԥ��p~FQ%z6X`�u�F%���5��jHT� '}lԮ�tyt��^�����䯹�R�\����NA�N�y5'e�D&�&p0����VU!Pv;uM
��Յ�K�H�\B��"�Yx��Gu�v���&c)4�KE�c<��K�Ϗ��B"ν�!���	��E�"�kccL�����)7���8��S���/x'M_e3���}�>ߠf<GC��f���ڑ39�xy�<�
d+�����S#ϔe&i���ȋr{#�:�����Z�TEdr�8�Qg��ri'~!qr��
������K�[u��h F���	�U��_�B��X����Wk-�`rW lPN�"�OX�=/$��%;8���
�s���݈o�����_���Y(�N�'�g� 
��Ә�D���Ð�-�]J�bٷ����L������r�����RO~��y>��仌��D+l�O�~�j(��&eR/�CF^���Ćo~��Y���u���-q~��%�	c�e���H$�U}����0���D9�N�
��+oV���f4H��^t��L�i���;�S1�G���wyQ�_u�i]e|��ǐ2���;2.�X����X�f~��pG�A�P[p&��Q��Plz'`PJ�������+ɬɒ#����@zTeC�t���b�i�\��Tۿpb��N�'��l��bGiϼi�J�!�6t�\�Ir-a	Vܹ�VDbÐqL��������0�w�u�h��h�%�k$���d[p���q��G�S|{}�`�PeN��gLfmL�{�Kч�Fã�[܊�*6�jh��-��n f�]1�&�v��Zp�p8ሰ\�����f	ľ���i$�[>�f�s��CRq�qdΫ���û�د��\@z���	�F[�T��Ix.�뢣b��*��Ȧ#��s ��S��)rTq�L�t�{�~�B梓��\h�/�Ɏ��6[n��7�
UR������9a�r�wo˚�'ѡ�­�s�����2H.���s9Cr)i�,p�.UH4����#��jAG��{�����l�A����{�b�1���k�+&i�t�3�)�7�����T"࿚���1?�U�>}ܨ�Ru�~��쟈f��j}E�bFR�T9�"�9�)wGNf��c��h�BN�e���jv�֏��	����*���0����2ԡ�6W@����>vgT�]�!S���VІ+�ĳ���:��7���g-@��� ��l�x�JI3B�#�*а���mR�����,��xM�MD,m��k?���Γ9-,���e��I����/nu:�?� P�����Չ��'�U|�+?iNJ���B04wJg��7����Yń���:��5�e��F4GBOKi�}�~q��·�3�d#��Vm��'ewY�P�[� �U�-�{7���5b��֝�f�wCXL��\�P����.���#x��`���ЖaB�-J��Ba!F��Op�L�k�y~M�@uT��$�Z&߼�N�4���d[����T�K��:H�����/�8�Gy��c雚�e]�8��^:�b�Ǝ��c�xQC
��kZ�,��k�����%�¾+���KFF�I�^��&d�s6��m��a�C���hfͶ ���k�Y�5$I]��ҷ�@��B�k$�	��$N�N�S�@
���	��1}R�|M)+NaZR��;�Q�}T]<m�����nJ|��>�i󠒧�k5?@���t#l�|FJ�O�>�ab�>���'央.��M�f �x=ryT�}�ů�1�䓚�<�����Ha�k�_;����.E9�"���}���,��G*Jv��7Փٰw�����瞱!�����y�fa�����l��_� �&C!3$v�i>��x�����P���T������6�@޺�@���kH 1D��B�G��:�J�ʢ��Xh�w�n��/���L��^��K���#�%�c��uyiD\d��B*	|�"ˏ�	H��yh6�gק_�;�����J�}�)�7�1�s�n���r�s2 faL�/�`�M9*���2��.8�p܅�HU��e5��=T� �C�p̴(�f���U�,<k��M���_��L��T�ٻX�#�PkԽ���Tzb�a��^��&w����Kx�E5����2D�Ӏ��B����� �tS�����`7C��]7/7@���-}�g#-ŢC�R�L����q�?mQ@���@��=�a�\�}d���5�\��T���I�c��������S��*�+�<��wy_�=�G�ǉ""�1����ML\<���8b������ˢ𛅕:WWv���iّBZy����t�x'�z�p���AP��(1��٫�5��M7nZ�
�Wao6m����	X�`�d�������*]H���&��E~[.+yKN��	ǌG����@�𐃂p����$/��ھ���j�3�X
9����s�w��
='����6fL^.1���aZ����8��tL��	��x"��c�.OT؇�E�qP���!ѴK�B���dL�j�t���cl�R͕���ȈTu�X�Ƈ�,��sw�H�[��K�\�Qa$xY��ƀ��$R-�����d�0g ���|1zV⿴�<��D���^]���0�D��������6�Y�����-�t�4�%�q��\`�ڡ?W`��|=��71�����8�{���՞�&YG��%/��Q>�	�;'8�:r�lЖO��l��w�{�;������� e�������F��!*%��������;@����".����zX$UEn9��Jz����P�h������Z���"Z�{�wm⴨x��͓'D�n��#��GP�q\ &�n�vL��cz۽rY����N7`/��o$͜�՞��t�z@�V�u*�^wk��$���D�{YX�i����Ȭ���5b=I;x9��%z%��}M���S��T�@Ձ7]������1���w�-�CE��5��ژ4����N7��U�+ ��������<��a~��'�h?���
b+%C��y�fJK����)�W?�]��S2�����v�a_d��s� L>҄Ot1�ۅ�LK�VS�K����s��-<i�I��%�x��5����j"d�:.�o�ú����	�#1��$B�RT?{�}n���4F���M}�RI���ź+=Ea����`y	�-�D�D��9��x�-M!n��?���-M��S�'���;��E4������B����7�7�����<��.D��D��f�3i�/����5�-��m���0Dq,Y��J���π�9����TDnӓ�,!Pz��y��T�)R�#ڲ�}�DO�$?(��-#]�g���ʏ�J�8l-�{CRĲ^�k��p��OpG��Q)�_��㚂��R"�Ŭ3�ՊPC3 ���RGG�q���CӴD����r��"?��[�Z�>M�~k�˭q��ooH���M���h����f=�����������D���*����9x���bV	�fx�w:��^�H�+�]P�0ן�=�3,�}9ɾj��<��[�U��R)#؁�T*�L��5\�hSL#0�v�zL�������W�s�X��Py�l�qU�$z2Pgs��O�^0�#���4���OPa?���
Q>���#Ë��
�'�x�I'I�ܐ��v�~'Ii�|�~ �@�qrK^�Sa�K��p�$��a��/�~�J�xD-z�jn����[�����]�<���/�4y�o�|ul�O٪�P��;�������ѵ�踗i��$.���ĝ�k�ʸ(j�N28���V7�&e�L`}��u@�x�荶�:�W��잡Ff�o楛��=z�q��φ�D-G�Ѥ��;��2�U��9d��b�����
��O���Ό����: H&����S���O�N��_�I��6�[� ڀ���zc�����W��e�ho�o��w��w͜�,%���u2�8��X-`K��'o)G�{�`�n��;DP����Ԯ��A��i���B�OD�}�n!G�akM�_�1�Lᅿ��|��K���T
�l%�G���x8:0"_�i�L�*j;휈9�Ɋ�����J^Mm�v
/��>����K���4xL�Bʁ�Bؙ�9��Ԃ�fNQ�1@NKWt�ϩ�.y�х<K���!}8�2�oS��4�࿄�|#�VP�������Zy�C&��Ę����KO*�<]���b�c�_s�_��7j�I�]�6B��J��7��46i��6j�<���Y-�Ȉ�s���������;Ҝ����缈�w�l_m��oN{uB�f����io�kxUU�-��O��R�a�� ��0��3�������O�g��@-i{DC�v�������WΘ������G��xʠ���r4s�;�;����f�<��P�A�����i�b�#��=�&@�1���-	,��Gp�3��Q^�=s�R4���7V�'^�R�:��<�R��w��o���ӗ3>�G��g7a�I�a��]����7̀��}s鋽����� /�a�;��zؙ�!�~7�5�s	^,�{G�+���@��O�⦆�ʉxe�#��;Z��3���Ii�����F��u?��!)�����<r�¤����?�*��zAJ�M}��v�g�a�J��IE%��ذ)��A��р,��~�E��ԑU���Zӟ�jۦ���Ӻ���5�I��=瀅O-U�Qm:���3�`'��+\�X�^�+���=�z�}�	��ɴ}pq+��I���8���h�39��asI��!.z��tU��ޫ�*?u�,�!�W��T��bF���pq�#xw�����9A>� 5	lrϛ�e-y�F�X��֯���\��~nw{�w������We"��j_��2n�8t���!��J��g���8mprM�E���7���`����Ӿ�fU���ej�xѰ�D�T���>��"W�v�qu�hs�H���*�y0q�;�D��~���U9�5�ҽ"�M[?LR�~�H*h	�] ���$�q3���L����$Q�^�ɻS�z�k�����������2ܧ�?��j�F���V_�W�))8��V+W!�����@��6�[��?�y�2�� sQL�B,��星ҩ$�"���H��v=��H�*f��Ct4�b�(�S�K����nb��WЗ�OB�����,Ju&�(��l��;wP�;���Z����ޓ@��BL����M�ԸCl�kXNV��3��b�6���IKa50/�x�a���ӫbj!5Q®���p+5*�������X)���D�-Dm
�����˵��wDG�Јz!
Q>��r\�{u��9��Df/�� ��ֆ&0S�ֺEm�B�6%Kp؊@aF�,.2p~'���t�����Ak��#�*F��w��G�1p���>�l�"�n��[W!(�m\D�ˍ��Q����@��LMɑ�|%��-�����\k���'�^��s��+[���7�:�(�zn�'�z�03�P:zK������5y�n@�8���>�h5�9��AE ԂC�@w��xp���^�o�r\�x�kC�k���垿��z��I�� œ��}�zc$
��n:���g� +�6��ܱK_�T��;i.�tk*��8��\������F���
v����vؿ��(�Y�7����^�3,�eTzH���,�b��2$L��g�Ta?���ewt����w�;08M�tB�l})U�s�I]S�X�{�<�j�����w~�|z�x]����[� ����D�Zo��
TZK>�ZRZ%��,+A%�#1''�D�<c��̧����8=�z#��K���	�QxT�ll2�ǽU�{._/�;r+��}��u���i�=��H��䶘D�f�+����k���&=�WH��4ϯJo��6.V�<��##��5���o_��$��k�L$�<�ZM�ǎ��T�F�a�Ϛ���K��_!�Uۗ�xxv�?�y~���Vl����b�A�b��c�+����;9����>mE���?D���{N�PPV�Ȇ�A`0,�|b|EH���InC�����z<2fO���r�#�Ωp�-�7������V��L7Q�(�:��J�Ztq�X�4����p4|(~K�x�HĀ��Y�E�v������?��1o�q�Ҭ�;���q�O�t"_��M�թ좃X;j}FC�nS�q�&�s�9�〖U� 뉡5�y8l�[	*�	\�Ϯ���[){��c�/t�8����%@�R��[<	0��Y��{�fC�:�d�$��m�9�D]
�3�h�I�����Dq�b�J�2�����8e�]�/�#��`EZ�Y�FCe�hE��B�|�j/�оa:�,������-'�����̋��D��b�J��^�H�%��n!*�;�aM�h�����j�b�޷�;T�v��u�;:�#�Pu����ǩ'Y�_��g�C�jR�r�PI�dy�뭾�Y��Tv��nE�Ѣ���!Q��xq������wX鿩t�[?E����5U�X^D4S9�gʝ��3�@Lz��(�5�RKх����I�
�C����թ�w���2��ٚI�j�&�~*|��Qql�L���S��l��� �%Q��e�r��Af�`���F�齗�X�ߘ٤�`OC�����cY��`�S{���%�qص*r�|���n����M����!j�5r9�����B���V;%EU�׶<��Z
_#v��{�}]'	q0������@�T*G�[^%}���Q�����䗹��uh�ߒ8�P20
r\������BJ��[�S=�ߑ&@��#���ar�ERN-35�M�GO6@�z��W�>�03���#�[���1��k��&�*ҹ�������l:��^��jLP�67�������Y�,t�Hx��*��<�\K����5-�_x��۳�Yf�7��C�ݔ�"��7��Eφ
�/j�`��iS�y� ��W؜0�L	�e�9���4+OE����>?׻�������UI)�(?�RT�04��O5](���k���+�Ӈ�&9P�R��+���_�7�M @LVd�:��`cvFH��-X�9�׸�w�����d�c�e._�����L�4/�����go�9�/O��e6�'�1��s�d����n?����S^"�v>��Д�J]!����?�)r�g#@1���cb2>x�;�.!��R�Y�o"w(���+%����:��� ��L��^bV��3e����l�JC�b��-�MG�d�{�V���'Һ��u�!ξ���ZTD�����/�o��C&�i�[N����7�m=�[��������]P��s��'a�����#;�;�'ޤ���ҩ�ַ&Y*4AR�I���۪�	X�J���3����C@�����In����l���C���	�܇��k���=�}�@�\��9����?|0,�h�-W��`d��^�Ǒ�h6��̙ �ڋz֦\:����e9�M��#� �z�;|��:���H�����\�('��y� 6M�7��(	Y�Q��Q��Da�A�~T..��eb<񚛦k��>�?*�J]C�e+�����$PH�#�O������f��%���̢=�ə%��+���o>�Y943*h3���3��k�����o�̜���5�hS�]�R<5{w7���^�hR�Q��׽s�RLT������Bǣ!�;�ۋ��������E�g_���|������ȡu9�Dd������`��[�����k���M�|G#�r���;d���[ߐ����9�m������z���V��<�'�	6ֲ�ͭ����)�uۇ�����E.����/�&x#T�kep��d1!��^��f�����@E�Ջ�(@��zY��J\��V��@D���́4x��b��Hֶ=��_�۵�ژ����kZ+��	��uUu�Jq߾�-����r�>��"��� �(�m}����z��X� 2�ʿ�!6[�;%� ©.�Ʒ$y~o���/�2?��On�սj%���t�˾��l^��ب�=�����ͻ�3s�4�~	��������(�����rb��>
l�0� uN2*�C%�4h�ջ䋼N j+��˳�D���%]��I����] �s�o䔷ZD���ƋM�9� "�a���y���w��᧛7�h?`���n"�AG�~sx������1Z�-��{�!i�P���'��V+���<=�>���K�ѱ��_��M;�T�PJ<������۹�=�{BÓ�f,�^���p��嗵����"�Z��ܮ��hU�.=�L~d��{p�k2#�/YRK�b�ˁ��9e`b���j��D���l�M��R�]�M��G{�8!e�C��������&�x�"q��a`]��i�g�,ՊfX-V����sg�9˼b�z��g�Y���O�l'͓s�,����n+|Z�A��M���p�+�H1�у�'-���_�j?��e�C6J�(s�6��+z# D�U��Ȳ:9��S1��9\5�':��à�s�X QN�A�M�67��βA�P]��4�D&ɍ��A0�u�N~�ä�eH/�@
Us�hh�$��&*�F�afh�[r2��9n�ϖ����Oī�N�Aj0X�cAmr^��쭇W�~�Pz0����^yM�f�@��XB�E4���w�{ք́83�߇�f�^����t�{�`�	O�@�i�����5�J�w���}���C(N����ت�� h��R6*ν̗��t��e��he	�zT Be`��p+LIP5��}ҧ�!��'�d�)j!8;��μM�1&f�ְ�9��v՘:�݂�����4���Pzb@z֑)��}�?51>�ƀ]CRK.�'_��C�35	�@��i?�kh�ł����nk"��ж\�~j�!��^�\��Os��GO4v�{�é�R%'B�u�V���4�9�M���������\վ\�0�/:��r�O�l1���i\#��\�
��B�8�r���'V���F�J��$9E*���QJ�jg�˕��K[#ܚNc�Y�A�֩r��~�&/�[�WqTN����ˍ}|�K����&��oȇ�	�i$��*�pg��a�
&�Bʀ6�h����J[Xy3b&�D�֊��P)}Zs5�SyG�%f���y�_���g�kh6�Єo�$u�_I��ɇ�z�r�!��֧?�˹nS�8��q�bźo�ah�H��$(}�Ѱ���$��Vv���:���ly8�)�R���������S�?W��4W��X�&z�H-����N��l{]��T05@$B�x���Ŵ�3���T.X=��iȔV�L.�Q�Ƈ��҃$���*�!�HO�4��D�����-��c�Gc�+'G�I�V���w���Rh�Jb���T=Y�W�5���A*K�`��lw?{�~�����s#^A��E���m��qg�����ݐ�o+׬ZGm�*����Ⱦ+ �\�+�ܼ�Q���p����>�9V�홵��d�%ek#AX�*��{�~.ޥ-�����P�����7��l�޴�W����m�\�	#U��h�ԥ��޸HE���S�a�?�� G@�GJ��T5S,q�M�JH���>���* �3W�噊ڋ�;���	���jGd��]\�����Bf�P���M����f��C��`V�n������x�A��Pʑ����/]�9Y緹����Q0�-�T�D�|9Yu�h�i_ C�yDmH��m^1���O�$��`�ʻ��G.�+E�J:3�SF�1�|6�)�kVBb	px�%Mte��{�@��3�q�u`��DY}ʶ�#�3��}�+]$�6'�� ��;��i�iNrP�Ȕ�RT�% 9ʧGZ0-�{�sX�(�����0�IP):��~��E��](�7U�
j���L:�
��i> i�m �#曧��<�v�l&�c����Z;�cv���ۣ��o�T�9�����h�G�?.�3c�[���Ԏ�əvZO��9rن�PyG7CH;�t�[�u�3C@����,����ԫ$/�h^��V��͵-�X�^�o�J�ɮe֎.������m�c����T�67\��^��!���n�� ɂ3��J�A�	\���E����c�W�!49�ٞ��)�=)�g�jm�kh>{=�T�S�(M�T�Bʱ���U>
7YB(��`wq?"Z	�����&F��ԇA��<q�,��/� �\�y#�Y/$���>�N�5�騾�d���^��с�ʲnɵt�7rRk�f��.�1���,��1��I��
�ƕuMp2���ݢ�p�FLGݭ��5���b��ͧ��p�O��B�/��U��}�U<��s�X�:�<��=�6�������"C'���(�GPU��`��4�Bs�U	�T7*v��ړOdH�l�'Ub�P?�})�U�������L����.�Z(	v�T%�7{��������<����x��v��n>4��OK2�<ƅK�h��;�+���"��f�f����QU��5#�ie =�X����V�X� �nD�K��
�#0��~fz�sFe�h��[5�8���ܭ��k��"��u�F���~BB�k�M����Qc�K���~�ƛ������K������iqUf��[�	ha�b��%CBw3]�!�-��S�������Q8G���U�@��'3��<lN�_�t�O�vI�X�~)q+����4����Z����|�^���;0#�SpB���UUAV�m�-�}Z�?r�����׳���a���"%�cZ���w�F>�&ٽ�̍�8�*T�`���ٚh������Q�
�O3u?Z�F&`V��S�Q���v� 浥�r�sg O$yX�d��Vko2�����Y0S�S>���u�<�����T�������2um4�Yl/��9M�����?�'IQ���z?]�uMJ�
��(AW`R�y����4z��UA(O�`<NUl$7�/u��b�M�Ei��D���T�n��X��v��V�.���e!%r���(^hr;�;�{�xz�l�[����hޤ����Nf�M�FyR��}#Ԇg|��f��B�wf��^���~�N�YY�hE�����Z�<���P8;�z��Lkϙf&����b���?
��s����?��N0R�_��%.�|��F���2�q������f��;��P�ɀX�W�^N��E$6��#V�x�K��6[�'8�c�.�"b3��-[}'VߐIp���&l�J�n��h��9�]�nA�{������9��N��w%?��J�4J����0��8R$f"�U�\G�i.���"t��[	��p��g��)E>2>J�~���������	h�`���
����J:�X^���~�XlxV64EB    dba2    22a0����$و�h�rhrT	=��!ic��_�[��G��-��B��֒�a�\֠�`�s�����؄�|T"=��
Q \�yDk
��*��ߓ�^�����<����[�� 	�P􅁋!�5��?�o����R��t�x��]e<�`�?uj�����a:e�9Hv��HU���&�>LRr��+�F2Dr9Q!ØV����L+��U?��%Q�PJ}Y(򤢓[3�r�W�e�{Q3gS���P|C��*�X'��_�IU�x�xq��|[N�Z��U����z�	�[��
��a�].~4���Ҁ��ab&ߢW����A�e柴qFG#�U�- �#m%�%���t���Ls�;^�� P�>�e]�I9?�֗�-Ih+�"Y櫡�
̓�9���{QR���*�)V��Ǩ��T�K��*���>ĸ��X¿Mj�D�\.����O���v�+�����Zn����nG�ҥ���2q-lh���&��٣}S���2�Ս�$-��ϫ��TY��*��+����T,gs{�?G�T�C���L���H���4^K�g9q�j9j)���cF�Q�1����H����&����ڢ���R��M|J>='@��Yv�I&S$�?�"x��;�p�DNS���)��~��qӡ��<�a�TfRS�@����c�1�ʩF��ZF�L��,b�}����I��*\pϮ�h�N�t,�U�ڊz���c�Ρ?՗&�K�v�����U�h�eh#"k��'��F�v���P�d�ӑo
�1�� �B
�$��u͹qP&l��ʣ�F�h�]	�������QG0��n}o,�[7�.�Ҿӹ��^X።�yK]_1�2B�
Ә�'t�dҡC"�?����ޖ��O�yF�a��aKHsk�A�[��ՎtR/J�N2������[�(�q�9.[Ǔ7n0�����5�ZJ��T������t�<�2߯��X)ӏ��6I�ZfW�=^&DI!�~����[`�r��ۉ�0~B��#�����	f�X�4��Q]}�?�S�F�$�n�g��:Aܢw '��6>/�������1�8<�^n' I�CDGJ�,c��Th-�*O6���������� �%��Q�(w1m��m$�8⠔pꠍ(1��#~�[�}H� =M��=D	s���7)�y%��n V�l���!�"[�M�~À��U�$�Τ����Hܥ��F�
��C�V
L &yN��;�L8�G�\�L��O�޼�C��ɚ�2��3y�bG�g�b�(wV�F���f
�l�q@�E�9�iPn�]s�$��lZ&Si��X��9L�2�R,�A���b�%U7����Dj>J&��eq�������b��2`�!{8���HE�n�����l��k(k��1T�1�+9�0VV��moʸ<�K�a�����g��l0{8V�
tUf��,��o��6$�'K>O�h���b��"�S�t�n�X}vq�m�d�99b,��V�A�a*ʫ1D��.Il���[-�����LJ�Ў~۟c�V`��iF`���q��%��,��E�Z�ō���cj��CG���w�8���Y���S� ���GLD���z\��{Ĝx¼��s&"ʚ5��
���.���S�7���[��5�޿��	��d�;����Pҫt���ޜ֞�-s�{"�e��PX�(����mGP&[��" ��<᪪x�ԣQ����+D�i3w[��}:o^�2�Xx��+jͽ.{-�k�ɬ�V�@	�
r��+��/��rPO��id2�h��%W]+yEv�����6�w-�3��5��l��V�Y�i�/�F?���aeZ�� q����6���#�~��}��˄c� �B]X�6玓�Å�`���;��7u�)���3��j�<����)��Mm[�������Ü�~\�t�yヤ0���޹�B&ll��N��4;��Utqb�9�F��#�LJ�����N ����3�
�6�4��7.8	��\� с)F@��xG�y�P���}�7�]�a�"��-��2*��ܩ�/�N 0�ߙl��h���I@+RGt��M���
�� <�Kț�(%p�������PyFo��|�3�?rgګ�8H#��&JgxY�W�B����H} ]�Z��A�v����P�c|^�a��<[�m���Κ���֨EU��z[��xeM��W�s�pN|{[_��@��%,rKS�»G��Y�
z�AQ��<�C�ԑ��{���;.+�G� �1�O��k��;O�j��Κ�g�7��TŻ��K���ѭ����zG���i�w�vh#�glEg	�!�c�IZ�D���up�� 0]MV�$��AcB/�q�%�k�����tlQ��w��م8�Z$���9��=if� ��@�K�1���I��Z0��*���ܳ��mV���Y� �3����-�w<��2J���ϻ�(�>dy8�ؼUT<��S@��o­�h_�}�Ë"U�h6;Bk��F��uhsɊ�1x��V�0�X�$C�4{�;�~n{K]9Ơ+�L�''�r?�-��@��#�W(o��q�B��(�����x�^���Ct�����sÑsma�R���kO��nH&��2,峰��>��q��v�ț�7/q�<��ע}�ҺQo�ś��0G�/O�ߟz��3���e�J��,AZ�F־�8O"`�87en�B��}��t3��U{R�¹�tph�U������ٳ��-���p����o�5�Aq7kĂ��q�e_/rڳ#vC*�k�O��`p ����Y�)�(Fq�N���ߢ��/�$�o�4lr��އ#��qpW<9[K6�"PS_����O��{�0��?�&��M��L��̵�B��:�� $;�QU��CA�L�?[-bI��4�\���2�>�nn��b����9�n+2�M��X���01�8#[{�	�8+:��+36T
$������
1�GEG:٢�j#��Ď-��%���I�$ף)o�<�;�ɡg �nx3�6�?�8DӕY(9�~�v0�B����U���j?oh��AW�[���`�*��ԅ}�\m��l�y�� |fBJ=[�i��#�fDMr�����\��7-���^\,B���%t�cړ�.!�bhK�,n��Y]�A�z�=��Y!_T9H.gV!m�� ���MG���jT"��κe�!Ց��S�h��͎�%c��~+�g������hZ��\h$2�`�m�]���*GZ1P�HHM2��E����6�)�C�ó�:-*��5,^K�+�֊ΓKg[WX���x��r@�r��82��D�{2��+}�'@�p`�kjK�,1�G\h����VQ7�pbN3S;ogZ.���k��G��B8�w��py%�u%���3��8ln#ry���=*D�ؠ$G8�O����yz^��z.M�Mc{YRE�K�/�p���H	5��-*�+�PU_��p�!����yo�\�L���	t�ihr��r�.�_���<��@R�t��h�����>4ʆ���&��u���sF�؃(�S��_���sEӧ[&!T�kQ�; @�t�b`H2&�����/��V�ݒe���'B�����="(�C����9�
����}�A�s�ǋ=��_@<��-��|#��m
����� ��s0�~	�]���:q��%#�Ө�H��`_���������@�g�̪��&]M���cZ���Т^q	��������oO�e����,|q7�3<2Pyz��4��m$7"X׫ؼ��(��=Զ
�ժ�
+�q�h-A5�~�G�$�?�l�ă�����E��3���Oiq'�<�V 3�w�Y�&�)�\e�?7��M��y#�Ǆ�+2��7b��@����b	h���M�в�Ϣ�j͉H���r��P#�ª/B��l�����H�ָ�
�@o�$+����EN;�A�`4�{u�8[�T�v�Lr��:1��h�Aԙa+`ߺ�?�V ���1^=f�ϠN��s訲Y84���Tƅ�TK����L}����T������ƺ�u��F���^���ޠ���.����V8~�����h]IA�����U�0��~<jg�դ���������p��4<>ޔ�?#J��L��TJ�oB����� ��jH�&����9SP"������;{m�RT3鿡B`%�����3w,�������w�S@q�4s�i��A�	�~`1�s���0�ݵ+>c�7􃻍���B��Lx4Q�'����R�R8���@��%j��pê�yoS��[}�vd�@k
|�����(:h�M�R�q���i��\�Eف@��N�;'C����Ag�PhϿ蝷�����޵Srڅv[]���"t.Q,+���iP�E����>/w[ ��2��kտM$�
�S+��+�jh(G�g��R���M��:�oa���&������?�n"Oq��s���kW��x�at��L(��!A�O� �W��s8�0D�J,��~<_�P���e���L��l�M3@�L�o��Ϋ�`84�D!�� ���f��wd7��M��[���! ���F��E��n��F��`g*	q �[q5��,�R������~��F@,	ϓB-g~w[m&�!��o�L��>��\���Xh��P�Q\½�\vP�:�GU1>���nݾ_p4=�	`��+�,�hT�Z��pF.�m��NZ5~
���^~#�e�P�\j<'ǔ�F���b���=���UP��Ǽ���ʪ��"�_,\��P]�ǫU�"9��u�y��!Q��P����D�JY�ƪ�Y����%�bfr���ݨAۑ�F��s'��.��&�@і�7847�XI\�j��xt(� ۇ_�K{��yWXoC���[-���Hw�F�f�o���y��N�V��T�@-I�T���N��z�@����b1�D�<F��}q�\N����u�����Ͱ\�e�sM>�v�B��@gG�/���]v�I3�.�n�͕�^��b���p�jny�����&�ׅ?M4X�����(����.���Gf��	�?=�d^��	�g�P������A�:7yɚ��{��(�%.����`;���H���e�j�yN�(�MwFy�������%`�Z�R�>��:��^ ���w]s�f��\܅��o6�6HA� ƭx�E�4$3)��@Y�-�b.�@�%�/�`���ij�EV�l^a�P�|,]ş��
|k���� aC7�ܰ��Z�YRg\ �	b��Zi�1��:Ɩ��W�gޭ�Iꍸ���^�Q̧���
	��X��_�Z¹k>�(��g��d!꼴�þ��c2Q"5m`�sY;-��@�]L��~|v��~թ�ɻ��Կi�0��k� 4-��u���t�J������G /�]I�_g�P�c3珌��ʽα�n.����~�qEs2�S15�$O>�^��M�#�6��`��A����<�,l�I
�>I�:�Ie?.�qH=����>�T���gɪ�*�R�|m���<LL�$��)͡nJǏ]�.S|��.���E؈��;F=Y(�u��Y�x�xμ}�6t��Vϟf��	#�<ۯ�j�L�BJ�W8/��2�>��%�_x���U&P��z4�L�Д73�л>7����2�u,I�N�û�'�j�[��e��G�ݎh+�ˮ-��z��tjL���%���Ȼ�@�|٤��Nxi�֖Fz1XYo_t�[�4#�5DN�uG	�����neӜ�B�Y�x�nƱ�ޑ~j^G����^N�?����/�*j�Ko7>�q��1����~���\N���?B:�M �Em-&S�c�K��%c���#|�Ÿb�Z�X��o��\�R��� �i��ϗɺm�θ��?%�L?v�ע��g�L�3ۇ'�?��쏅��X��|��K�tT��@�.��O��_-�,I����U�t׶�f� v�~G�x2��/2��!�bs�5)�q���w��#�S�(���ى�-��@�p�'���.�ٚs=�8%�g��`�=�v?���mg/Ҏ5���R@��G>-��b� �`Ƃ<�d����?��eZ_��KVs��pPpA!�GPQ��r�&�4@T����@m�K��;�/��pU�iH������3���0�y@�a���3��>���K�1�G6���^�(]�l��X�����ؽ�.��χf��/"�T�"�UQ{+�QN�����e�+ѩ}�X��&	*!#J �� Îj0��+���r��g�P3s��8ɿi�:�������|>��b0�54����Pѽ�d ��SS�F�oȑ�vc��#�}g��c�	tc�O΂S�o���l�%��	z���I#9��a|zyhg�ҜG�6�BӾ�/*2F�L�B�ji��؝V�?)�%�5��/�k ���eP��>8����
�$��Z��;����%�;t�s/���Nf��@u\:�?)�A<�g���[l	�u���n5b��hv���pֺ��b�	�g�6�A�Awg�f��3a�n�o�Ӫ�\)QɊ�%>	�g�b2�=��t����ȉ�]0Z{R�m�Éx�����!3�o��5���;����$ƔXR!�p�	� -s�,k5��*2�rކ��<vC�����vЌsҒй#��X�s3F"��c4{�Bǈ*�cc\��lX�7\�l��d:��f�$��[��6���[B}���g��?�����m+z�?�KS��.��@�NGɖ�s�>}��&A��u��wBqvT�o-?@N�o:�8��i�:�e��HQ���M+�����/ �^�R�펉@$~�ƙ-�V���m�B	&�l��c���2����k�q��O�f|��������%uo6�F�Mp�!���m�>��'?��5{PKZ�1�9�fzW�/n"Ҫ��Ձ��A���]؟�
eM�-����A��4?�~�r1 ���e�Ź��¾�殾V���H��y�^�V�꼖 �4�O@�[���,����p)��|^�#�n�[�z�^��{��Z���3���RY!��X:J���Ă�ڳ�Y!�BQ�Z1��&�r�
[��f�����M��5�-a��B��[�Yy�w��.����Gɏ��v�����mF�|��AI��=��A�y����%"����L��V�҈H@�g.��+�%�`0����B��e�7}���y������E犸�S}ZL{�'*�ۿ����Jh�w2�8FЅ��&}�*�H��]������.�q�|��m�8$U�+*.�;���l�3�����nt,]]'���$�M�Pw�
)���ѱ���R<.� ��@e[�WK?�� A e+0J�ۏs�r�㸰�"}�RL��+������5�ς���rH7ɦ׵��Ņ��e�I�E����IoRؓ���u���s�}�P�O+�n7@�0Y�o�,�#�M�����qR���}�V�4!����Z8&��U:w��	�&�Wh���4��e��>=FWL<m�=B�3{ʇ�oO΁a�P��.������ }T�H���([v0��_�C�̢�[5}�x�lFO��MB�|���O�p!Ѩ����ElNKD��[��t�2�A��рHF��L�%��S�x.����u7�E���n�����d��[ۣ:�O��r"���:v�f����p��Y:1��csg�<��+&�R���2�7�,���â��`c�����e8�(^Q����.���G1�E�B�Fw,n%�s�,�����w�9A8��SĊ-�QP`ͩ>M���f��3Q����΁Eݞ2���"�:�.|p���C�GE&��D��8`/X�Ƨͳr3�}^��D9�����W��E�y�e��`�~����2آu�*���@��ܝA1	�w_��h|l$x��9��)b@u1{@F;�����#��A;Q_K�ϟ��JBA=a �4��(���J,�Yt(���v��{Y"������"%��8/��z6�OL�m6��Rg��b�iU�ͺy�J�~���T#cX@f��5�4�lJ�XA<��J�Ann���������8��&�k]!�d�isTX�Kt�U�b�K�ŵ����'�J�(��&X�m�N;:���X�@3)��J��ܪ쁷g�� ������ҁi�C"�����m�>�	�b6eK�ܭ�Z�!4�ռk:G'Q�K��6ǃ(����׮*�0bEv٠YAqz{^{w.�7�r���x���4@�����ؘj�� ��H�_I�0з=TZ�@B��!�`Ȉ��i����D�׆,=K��xw�E�}T�j7+��=�R��{X��G )�ؤ�j7Cd-'+o��3�PT%Z���p�ߚ�Yo�W3�?E�Ye�e�P�Z΂��Y+zN���}Z� �%ױIaφ��4����d�R�joH6�u�8���zь��Ɠ���]5~v�l���Q��RS��bψ��#�� W��5R12�n��)�i5/srF���j�A� u�*[�|\y��Bb���$�[�R6�:
�^��Cp\��,�(7��΀����k�N����A���u�S(s�!X����R4UqJ�eI3��pSm��������Kn��m4��Cɤf�����W�d�Y�������ѥ�9c�.�ݍ89Gn�)q`��O�?��9����B=