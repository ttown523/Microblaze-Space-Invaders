XlxV64EB    1870     6702svX�u)F�>�E���°/���X�]��\���}�l�Z3�:�j�Β'!�>aO��,�5Z'cC}�U���޷�O�;J�
�i�(�3^���`)� ��-��O��M
V���z��3��U2�/�N�[T����0���w�e��Sa��[�����cII�#�E�R�JdiD8L���� �u��E_*�ft+aȊn}�T�(�>�����`:`�^~�Dn��wj����A�w&�9EN�]#}^�T���f���!�x��$���Z�[��`I�w���VNv���B�-ƈ�c9�pZ"�a߂GY]�U� �?�[��!2T�O�0.�r�Jm9>���v<l�;�m�H�t%��7�PB�=N53�g�	s����{�̚�4�ڳr껉 Rv�ڭђ��&t^S�(')���H��Ί�p2�yPV�^9��\�x-ѱrPs9�b�JԤ�%&�2%Q��z���o�x�ۧ�b��p	A�KR[79ghl͒�ڟ�X+&�T�+�9F���`7���آY�3G�L����n:A׎W��H�"bʪX+S�7w�F��na�B=���Àq")�7��X�8�*�h�;S�Q4����/J �,�Q�,��2`.KP�ȳ/!~N�(�V�$0� ���OK8�+I=%�4z�o�x��(MQL��A�V����%�̢^�~jTIO\rw��/�d4��P�S��B(�B�����\�MS|�l[���^k<)��MG1�R�j4d��� ��C�y�Δ�VTA�(>�5��f��ڳ�8A��ԃ5��3d�5u�Ѥ|�_T=�S���9Eg�d�zhK����}��h��Ƥ�z�v�KP��
�h�,��zT�p�+�B�+�9�m�w�a�!��X�u�̢�'�T�Y|�=P17���u�|1�� �@��=
$
�:�BM��d�D��lmZ�~#Kr(%m4I;�&|�ϼ
H#�����nT6꼥9�sxc����v��	��U@5�	.?��1T�ß@�:�
�*!_�xx5zMh���{8	��!^�)Hv������x&A2a
�#�V�ϙ�I���G��u��Q�F1���k�y�t&�0+��"�D�1��_v/r�8�yϼI)!���nֲx[�tI\Q��1h<��/���PƉUV�?�m�R�G��a(�j�x. +�Z��yC%גW@�Ӿ+���|��^E��0v081�q���|�V-+]U�s�*B�J�J���>��������0^ND	/����%_@j������3v��O����(8~Tr�t������k.}Ԭ$� �>��>��e�a���0� ��d�l叫K�Lx���CLA��K
8�MR=�����q�XqK#>�m��0�a��${�hc�s�
�te<�t�xE#(;�k�<!���]�F�Hw`��&��_˒2M�ΐlW7!�
�|*�^W!��ի���B�\%⯃wqź�	�s�� jG��P;�D�o�jٙ^��L<}���PHC�H��V�}o�lnܮ�M�0���S�qN�7m����vD���� ցy��� `˷c阋9��2&�k�lSh<v;j�ٷ܅�ߖa��؏?f��3�]��<�J��;��p����E����o����B�sV1#�V}�Ra�$E