XlxV64EB    3bb3     f40�aa�$�Q-aV����4�-T�V.Ts� ?=����hd�f o/���r��C7gYD�궟�z�vjU�Y��#�;1��`�w�G����������Q�/J�5U��5H��7(��)Y�@ub�2aY�\��	�o���0"����V�c�����)�S�{��ad\�X3 ����08W"�h��O*c�����9~�㞷ƹ1�cxe�	*l��C'��3cڛ��GC�~Mu�<�b�C��������:"4 C���o�)����8��F���`^<ɭ%��q�ے��u�묶�ÁA0��81������u�� ��<[S 3to<�ŗ҅�7��CFDl��嫆���1gD2�w�~~(�Id �=l���Z1d-��QK�i	yW���)^Zdq8��]�e���P<��%Ƿ����]�k����.�|���Ο��(+B��P+��g��A���d� $���j����o��<;�����I%��q�B�J���UNxT��:ȂR)o�J�3�#���K?�)S�J �����S�ɑB�Z�I$���3I>q-%�[YEK�Q�n���F��E;]bUr#)�_�/��.,՚��y�� 67�=,^�Z�槆�c4���䰎�V�#ɔջ������O$����\SkU�7V1۩��F�������X�����!�/]����Q�jq`���S؆�Pq�\
�u��Ih����n�4�
�x9n�^!�Ht�84o�}r�B�(ɯ0����W��&���tKp6t^C�}���������7qr�qc���!�v�:Y ��\���[�a�a�*�#E�Z��vׂ���wzJ[{����XY���,�we�Kb�C�,UI|]��4����*��un������1�c�;��I�3I��~�y=�dUy��!���#;���Qڔ��8y�Vg�I�	�����3��^Iz�ЀK��ft(��%��ѫ3m���$"�m�ퟮ�ɓj����l�T)�Ғ]*o�
��0������:��x�VI�6����c!ٗ�YS����{�]�����MD��u�M�WD��޽���>��Ө+�<�ͪ���iK�|��;�d��V*�f)FB�*�d��=aPV#�q���F�2'��sJ�L#z��D�ؠ�9�����Ӊil����W��k܇pn���'*��+��:� T�^N�l*�J���'|�4��`𥌋(������#�&��a$��pDӭ��	��hd-à	�$I��A���~/�#����|�N��o��}Ā��\���Y��uQ~^�'�5c��;mj.��aU�w��v��M�]�Pf���Е'�HՓ\�:n|2#D_�i�
<�vK)"����A\_�='wt�x܅�
��OÜr�W�Kj�r���'�Y2�H<�Rᷙ�'+���h��j4�;�a��4p:�����4s�7��g��gM��d�x؎i֪��I��I��?MGJ��|f��
�1{��+���[�֚��L��p�jT�*�q(��=>��Z�� U1�ߊ��7@��:u^�C%8G��q2)���A��y*�d�eg���l��e���?�^,�4�hBT�?�шȅn�Cz�b'�2�|?(1ќ�AcaլP�+X`$� &|ȗ�4�?9�P���B����
lw��`���\��>U�\�G����e5R���JhRq^����vY3>���Z�?�s缏`,�5Ԣ���69��Ue�,{W�`�SH;�iϴT�ƍq���B��m�2�dB�:tU�OCT�ȓ3��e"-��54��I3�-E�>ʚ���H3����J|�$k�H\�6HN�>�b��Q*_T�����$R��\it)���1��
	���!�VH���{y6�)���R�tr�fV�6�W-�1�m�A��
7��gD��a�Cif�=�J��Ls,���(������6��a3�-s�h��;�<3��j����Z����j�2�u~��sk|p�ZI��ܸ��E��8�p"�v !x^A/��B̞��I��QI�3WE����*�s��/Љ!/�5]��a�KO��W/e]G��7�f�J�YL>�`8��ߎn�Z�QG��r�4w����8�*�1u��X*��MR��/�3�71��tlr�c�M�	��a���b��9�P ]@ʛ�>q�dg��8@���݂7��Eڰ�9��H��sA�����k�������ҏ�mZ����g5ȣ4����������HQ(o���(�1Ǌ
�=D������;;�S:i�N���T��"w(V�Ev��wT�B^]-����O*JG:��f��$}.��R�<�`�l���j~��;��I*��^k��Yj����������$CN?4�_Y�_�lWa�ذ�ͨ�G�+��8D/��!S� {�#a��̑]ĕ�59R�q�� ����*�'�g��#,7�R(�%�uQԤ�&����%�ï$;l���uV�o�7`qꊱ��T@�I%BoJhtp67R�]�-�+���j~�Ӡ]���S��v"��ѭ������rRF��JxP�j$_�ʒ�G��E��o��|U2�$��(ժ2a�ߞ�~5[=5��;&w��^�\w̓_Զ��8Y���m��Y��C7�cd���$�Odu�DqNl߳`�UT|�]�k�@�CIܙ<竘
dX�yԩ��܉�����XP��7�Qy�Gux,�Vt��iP���椚ġ x�@�c�ཧe��Gb��U�̃A�(G��B�O�NgJ=`�a O�j�p8"����0�8Ù������� _���h�8݌aX�2v7/Ǉ����0�ԏ�}�7G�Z�U2�I�%�e�ά�Z���J��p�9���Kw�R����J����������~�(2*2?�P�⮬�t$�_��6-����w�D�������P���^-:ǆD�q������9�!�p-[N�;:�SEWR��� -���2��Ǧ�`Ȍր�K����̘Q���0�j�LTE�0�}ּ=�|�g��*�����)8�$�����:cz���ԙ]�m�Gz7��՘��I������R����i������mޜ�X 
�}��,��T��x���A|,X�f�e���6&�mrܱ��<q�4g���j����2�H0K��v�S�&�����n�������`p��W���Ӗ�Oq�օ_�뱔�L�l,�.D<�Ө�˺f4����g�'�#ӄ�kK�O]�WA�1H�'� ��ej�oWO��:5'<7��%፥8ϽbH, ������P�'��X��Ϊ9:�%И%�i0�2?���F��^��cU�W�bF̂[�8\���/��y�A����,���w�1\o���=�\TvO��P�.�H����H����칩գ7$���o�	���<�mP���z�k��P�!���<*��p�1��L)����HQG̞Jyv���(�f.f����ֶ|��t�t}�[��P�a�י��g\�Z����1@T�ϧޖ8]i��Sm�,S=���#�/�t$����MUK�0��x��yG�� >��>�R̋v�SJ6 ���켵�1|��a饔�
���_ʯ���s�L���PSat�Y����0s�1V�5Q�u�F3v��5X"����J�Ⱦ �Bb��w��>u�m
KV�aB����zք�+��4v#���1`!L6m��� ��S
��ތ���D]�8�k��:Z����4<��#��-<�y'��]�]��:��u/:���Fp�� �ʾbQʵ�b��-��$���'�&����A��"|�8�O�W��K��ѕ_E�������C��l:S�.#*�J �ށ��y=