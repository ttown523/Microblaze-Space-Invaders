XlxV64EB    3f2a     fd0 ����Z}����n�͋mk#KÒb(tf�^*P��,7\_d�v��@9@����c��G��o�*��J93<�#J�O��o���D	�:!�ʯ��|�ר619�4���/�j�Q����&�S�DV�\��q�O�C�g�cph����*��@Í��{%��~��{\�B��%�'�M{vD�U�:�$��-���^�κX��>�s^M�/?�[����%2.�o+O�z�����/[#ID"���	ؗ���Cy�X'�It}�hحB<��B�F��D���\��?z��m��槪Si��Oz�}��'_���n9>����۪,v|0�L"���A{G�a�Yt񾆀,�5U��k��~S%ǘP��?����V��
�J��q��s��e�Z������5�!]/�}����"&�2�Wpr���1O˒�p�'I&QY��o��0;RT��y���4�D>d�%|�H�x"��5��b���1?s��xU�Z6)�c�"#_��Vjڋ>8�8'M�E���t��}�.�̵��T�/RB��o_!ٲQ�?��K�;���Ꮥ��޻I _s� >�l_�KP�γ��I��f�h2e���{����H=^���g��
B`�� c\�"D�+N���%���*���B�47z�P���Uȶ�t��O�(W��y���\\Q1x�����������X�g !.�	w�
���-�`�&-.�.�-�m�x�jL�޼>A���v�$Diߥ8DKsV�A2�H�L\4IQ!�85��3HC���C��`h�e���L:xh�%����t�5�&:�F�r9_��m27(jV�,{�ۆ
�Z���r��$A�#��[�r� �s ����+�� "p��w���lV��g�p�܊��Uub��|��V�7<���Q K���R #p���28�j3� ��+��D���K�3�=�`�tQ�Q�u����~��X����7 ^�,t.�\��i�=�Կ�*�^%&�����e���2�̀P�T�BB�n���G�DiO1�0�"V^�8?n�wsW�'?[�)X�^����Ϲ}�:�`%��	$�g��>ږ �Ó~�*��(�X>:pbѾ�H� ��$�s����^���E>�vK2a�UA�������p��>�6٣U���8��_���ͮz��<sS^�t���V��/w�3�PQH9 ]d�^b���	|��I
<�A�H��C�N���]v+�Q�=�[[�X\<���m�uy}�S� P�ɻI����n}W��?�Hw��]��Բ�PEɿ��y�y�x�"1h=,.����Zd���S'�[�$�f�f�2DE�����k�2v�@�_��'?���o��KS�"�� �==v4������&ś��_tː�&�I�[̠�p��A��,�a$f��h��QI�(59�#�y�:���EĊY�m�4l�¢G�yH`�Ok�CX��}�db���@�,̼֡=r�d�LD��WS:t�\���Z�(�yf�5�o�_��Ë���@�e��6�������Li�3���Ȣ�-��q1I��kԸM�а�g܋H��`@�v��;�w�	I�����ԥ�'	��Ƙݲ�|�:}T�B�\
30`�j���N"ZE�Pb`D�y�u�yԝ�Va}�J��q�m�f�Bfd�5Κ��8(D����F/���ƘgХt}|p$HV(��:��Eh�H����sD�����KIy����M�p��t-�e�ru��Ik��hge�+�� �K�gg]:�\�k8�ŅX�jb[ 4�}�c����R�3�b}M�|OoEw�֥���t��|�2J�9Wd���jɖ���b�[7gU�F�V�?�V����Za��	c|>@��ʑ�l��L��.�up���Ү��pP�@��a>�7kk�/�v��8Ƌ��`�ة�����V
7��=&*V���)��J}N�E���?�=�F�k�Q�c��0�&�����d��/���y�4	ӭ"�t���D���w�Z�^m{��N���K���l;/{���[�|. 6��&w*elٶ�VS��4����QmDBi���o"�9+�cu���P9!�}W�J6��D 0Q��\:_3Q�]|�������o�Gf�r�-�!�S�D����;�X�&��5�x�Ż��HØǯ=�f�d��:�2�*���,PL̺��v�C�y���9����6���{A��uv��PȬ�0l�܂�؁��06��[H��Iq�ÉApy����s��g��-�W���F���0��j����,5��Bc-���v��\�Z�k���է���Ͱ����%tn�:e�FE)������ϩg�@�e�P�|�z$�,}�TB!f=m�?Ud��!v�|��Qm�`�����U�i��61���]a�?��P�1�"~�)�����p8���5pũ՚B�0���Ae9^o�6B��[�M�fp['�Ť�h8ao��0��ɧ�\7Y��.z
��Qd"@����+�ߣ�����hݨ���OG�{���->�W8��/+��2)���K[��M\/�?�=�ݏ�f +��Ŧg-�g"����%g;�ڃ1$�l���nr��5-p�e����.�]�1�ӤQg�	�j=rV���7�a�]�U��w��h��*��aj�[	�u5չ�����]B	�R��������Ԏ��?���e��*A��)c�H�s��0Sy�c[m�������ݒ��ٙ4�p�s��82�Uo���eiP)q?X��A0���!LhL�.��krk��d��^��+����8�����˞������r̜ܲ:���aQ�[��z��/bx��򡇹��nG�GJ�9��[��!��|�v,��u��b�<�"��m3%,�J7mo�Eb��P�T�.gs��k��PC�#�{M]�o%s���,r%@<�"��6Í��ʳ>��osw�.Y��P�!��0T��g1����EG%$��+b*1�P���L�WW/X*���|W���sg�NsC�8I\���0n����.��B��Yz��`�YX �X��{�87�vc㗺r6*8_�� +2�0x�~��.���A�$k=�Q�ϒX�?TvBr��
��B��q�f�����ᗝ~x]q�o���t�ܩ��,Y-l��6�1�K��v�~G��n�Vna0H��u��>��~!�,�Wa&���"��'3��3�jν���0o4T	1��kJ��6<P�g`=O2�����b�)�$�S7�f����v�:�ag��E���ФKU�l��_�5v(�+���!ݎ�a��\7�d�����? ��@�c߬}�m��?�|��(�Yi3ޛ��IU0"�����Q�Y���h�en�����(�ճ-zP����sV`z���N�e�a��!��mHԞ�D۷�[8eΘ���b��D׾~�B���X��'�N���gR���]|��O�i��f�`�0�"������|�IA�ݓ'Z������P�@cۨ���{"R#�F��Ц^�>l�@���m�RW
�` �y]��6��W�;��A��Du�G��g�R���y��7u�!���~e�a�a��0g9>�bO��K��E49����&�j��.�6+���*�2�|���v����I�-ʄ�D��~dM*���B��u�S��~23��`�����XӏA��ta���[�p�^��ћ>�Nh!��H�47?yun�����Y���VH���հ��ݶ�fiߌt=���!��x�b��EA�����[��<A�d<a&���5YotP�_i%�b��ؤo�n��j�bK�Bq��
�������Ԏ������>���Ǒ��ѝ�fWYX��K@A^�G�a�V<�3�i�؜�<�(թ�����'�>bJ���{�+��Xm3��M �n	|���fN���r�$5f�����J����%4!���;��RM�*M����_		Rl�³�w�%Ԅhw-Gf��F�WE��Ո