XlxV64EB    2837     cd0�P�� �W���At�@Ņ�7��q����'E-��G���2�B��fR�����c-e��n�������h@_��~�W�n��{��ƯǗ�򏀷i_�`�d��^܍뙨�S�ˣ>6�T҃I�c�\��v�ck5;)*B���pwв��:m��
�_�$A ����p�G���z5�S�RDQV�O��:��gT⤔���8Wg>�iQd�:5�d&;��K��\oC7���Sg��A�Ȝ����	*<˘pr�~R��<5gZJ�WJYF��e��H%���Q�0/o�h����)�E9W��S�I�Ŏ�T0O�R>L�w�/��&j�T�K8E�5`��{ ��^�F(����u���2��s��U.[I�Mn��p)j�z�,a�C��]8 ��7x)��溴���pA�_"�~O�4g˯F2�v�!���?�����؅c஛��5��$�[�iv���4�ٱS@i�Lw���H���5<��r�->9ļ�QmG.�L��b��a�̌�е4�������3�X�n� P�%H�	p�?���l�T���^?-@���L�(۰x  �<�N���ִ�>�ʩ�I�Q�
L�X ������#��$j����*c'X_)/4��,�p�C�)~M=���Q?����r'QXEp��i�"�T�(�L��
	��y���:@7�Z��R�� ��[�"��҅s��mB��_��=�!ޘ��H��F9W�Ѽ
���Is�ь�T�M�Wܹ�_c�s���I���o����թ���
}�i�q��{�䌜�H�x�5���ms#!�7p��}&	P�!^�36�����~�\K��ё	�*��l�r��E~������O$���0�L\E�+މ�f�2�z�L{%8��4�D.�!ƭ�Њ�����m�
!11o)�����P��{�.���r;泺�x���8����-�D
H�2�k���b�I��Q�TX�v��@gC $�\ؽrv$��|��f�F���?��<M�w�J%�n2|��X^ƨ�ݎV��K�dpd��FS�~J����DW'��R�2�������L��g���������$TMX��~J�. �5pH#+ʶ� d�1Ξ `t�~~W��{=��d�/А_�j_fu�����4�OW]י������O���Q�nT�i�U�'�����)��N��uO��h��ø�Q-Ќ�	ZmD�[��������°���w��b<ًПG4_UռC�J����H9��2%#�w�`�r���.�GT,=�%R|��Y��F�!��LƓ&WT���/X�����|�q.����.[0f͍�/㞍q��s�]x"�b���#A~rk%i"{ �N����J;e\��w��{!�G��w5ф	��"jٴZ_ʝ�%�I���[�{��d���罵㚀3�k�g�}?����;4Q��{|:MsEWAܲ������g`R���a\����E�2�h�җg�ܕ;��ř���
�@����#��抉���F��ͬY���Q�Έ�4���=�z�$�@����.�8��C-��Be�"'����<7<�ި|j%��� IZ�^wd�fn�+|N��d��ib ��,;�咯o:��p�s��n�:���EArPD0Z�Ɩ�a��`f�Uȝy0@.�;�O.��j$E�ۘ�����!�"�g��e��*���ޒ�e�:,F|2��@�9'P���W��:?Eqn'/����_�Z�ؿ�
r���!;7�s6/�E�dA[���`��K罬}�$����+ߡ8;�����Ɏg��lQ|{���);���Q8�?n�e�YoQ�f��9��̢V|�lf��(�Y�C���j��%�X�o�'���E-�V�g��#���0���,�Ԅ�X"�-�,�:�Ŋ�2�Ʌ�_�8@ؐ��h�妦��<�QKI|]֒Sr3�dV�K ��y����+�t�S�x�9�x 2dR�"�N�ڪ�r��M]���*��%B��&b���M~�rbzg����'R�����gv7������v�\L8��t���Wݒ:�w+l��fsY^F�y��ѝL�c���H�9'�QcJ��ו�[��J�TKŢ�Tx@=�#�b�6��w�]�>�@�@Ư�U�㝸���h��%�9ٻ	J���w��uG�N����d[2v�'�v[jާ�����@+�\�[db˕�\i�W�j"���'ka��|o-qjY�8�fL�N,��D�	���#i@J�G<y�vi�s���5Џ�����o`��{Y�`/���L��!��H�z|��ȸ���2�g��U귇*����i'��sm����캵Vj:��7=�����,6 D�sJk��MлO��8�*.Y9�ˉ��%2I>���DA%�-��!�������AjK���)k� ��Sz��8^P��~O�x��xz��M���h��%\]A�Ԋq>24�����+>�8cC���7輪ځ;����#sx���
\��ʖ�8e<������gF�PZ��٤(\2��e߆��w|k��#�@�ݡәO���C~�{�=$*�b	1�N�Ti�'�$�gP��)U���Y[�����a��ȿu����d=;ݎ䌪�
�ɣZ�i��$i��?#Ki�N\:�^���E�k,x�H���(
��/7A�||@UB�myp7����S����X�?X��f&�������{�/Y���E�[�uc}Y��v�/r3(����pJ�7�w �	�KhNf�:L&w��+�Kp�\���l@�)�ٗm���
z��ؿW��<ɭ�%�ZXy28�/K�ӌa<\�X����~���QkW�(	(se��00��ʄ�eW�oy��maauL�Іu�,��-�;����<��;�(_ػ^�҅q1��	l*33R���1����_X.�JU�VI���e<�ՀD��Plk��ʿ��`��[�J�u���
n9��}����M+���%CA��Q�XDZ�}_�`��t�U��ҹã;p9�@�T("�ml�~ĺ�!���y�1OO���%�@9�����@14J�Iת���	�7$�ٿ�^����7φ����Ź��_��ʂ��� �c�/h[�ܩ�E�V� �C�&���L�9`eSFNhR��ƶ^�Ɉޢdi�R"��0��9�>��cz7n�x۵��s�2�����(v�4\�]��[�.%�2�=4jF�u�`��C�9�F�O�$yi�X?&j.�>���O�B����