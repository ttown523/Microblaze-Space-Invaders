XlxV64EB    4bc9    1460�>� ������ƖcL�d��l}�Ł�3:���`(�|U<�y��@n�Ƅm�!����̋��`a!��1Եm��+S�WU	Q�ҫ�l��*��&�ݏ�z��L��tj}M��*�_�B����|D������*/�5�%�����X
� nF�nd%��joy"sO0`2�F���>o��H�. �$ǵ�����(���/*�ڲ�u�D��k�>!�5E�@�I�펴�]CT��R_	M��;���,�@,�2����CpW�g���J5�-���?�a����/�̐7�0��z��C(�+�m���9S4՛J^�ѳC�wà��Obm�����[�,��2H�v���!nlJw{�
)S��;��d�*E�1��r����F&r��5�Y�(�����t���!�k�MC�̝�=�sd����E7�n��u�'Z��@�F���OB����x�[��>S�rC�[�4ػ �"N��o� ��Ր����:q��LG���N��Գ���@����(�-�z	Ř��`K��04�>��s8R�����`G%�L�@�@ǒ�ˌ��^O�K��t6-տ5����t $w̑M�@S���V��6������yW���.�w��+~��"�Ql�m�ud�W��2,f߶��V�$ݰ�\\;�T&�mDΊ�����ZT��gZj(�C��l	�I��}���6�
�k�^�3��to���*��^[A��"���X@XD�h�G�=��5��?΄u3����D]���H����cbPPn7b��e �'_j���=�rSuq��!䎒�b�pG@��3>R*�X�٥�#��f����;�-�R��>R&�Q����_,&�"��'p�A��C�I'��a�����ػ�����k|%����8�&�b�Њ}�u�Z�p��O��`,b���+3n^�y����}��[�@_�c��1+&~�Io�|���:���/���}e�%���$
g���>�}V~#k���S�#N�$#]��A^1Л��$s��rYdU!ϑ��1,5ux��[�οBg����5i�D�6�'T��iUg���G��b%�I����o��׼ѡ����	���܋��(�p���ʂW�x�羽�|��MC�� �!jd#���t��ĵ
M�^EV�/�_z���Ùm�tQHT ���eީ��~ة�<]$M�P�;�8g91�x ť�: �a�F�X���<��uB�Py��ΒpTͺ>T=��6Ie� �J�{�ݷBA�;���P"�P�{;`��|ƫuG�Pq����|�&��D�ÖB��K���S�K������Wx {�1SU��*E
pd��%��q'��rA�X�ᓄ�p�ro����{y��(�Ü� �B5���8��͊�f�S�Bh�?�E���{�M��ut&,j ����_lm�d�.v(]�Vu��2�����)ܐʈ�݊#h�;�i<��d�t�v����)�����/-��
���$Z�Q���o�o/�+U4]�H���CY��؂H���j�s�8��5˃A���Y~��X1F�|�L��&�4~d;�cHx���&$�"=��P��^f7jX�{�6���BM��IK��g���B2N���$��P�@�Ʋ%�,�x֨j)��H@��w��U�I�0|��o�����L�,9��O =Z-I�#(�nHc|,BÆ��rQ��v(1}�C'���l	y'B�X�?|E/V�\�*�M�0I�vC�-�7ƽ���~���5�oZyB�#ӽ���M���&	 �/���!�ߝN�������6hx�	�I^��L��0R�&J�G(0�\=nN��Wկ���3�j�q*Vjv��X�>5�����Z��i�em�@z)����i��Z7�өU~�j4�����?ɘ4weiG�ȉ��Cpa���6��T�9	*����_��)��D�n�}M]p�w�b�$0\����6�]��c7Kn��8��6��������6�?�7qE�TV��}�����iqސ-A��o�y���;�k��T"8˺�]I�{�%(B�¶��c�Rc��P����D~T�Z7�+|^7��&_6�a�ǃ��ym!o����_T�o�����iI,��k��B��2�aI��M,G����7�j�*w�?*re���Qi��_� �x���&��Z^���x��9�(�,m1�*wc�m�80gl��k�㢑"=�*$��8
��W�p�i��>�h�������8��^����B[I���w��h�hٜ�J�!+1�s��v��Z��߂�H8�Imϛ��`'b��/ ���(��&(2	R���Q��^s��\��L"|�j-����%����}��0�[�{�x#u����"���K�qN|c�p�(�M��|E;�ymN?��-Ѓ�3{L�M�P�Ul�1�7�;7<�?Fo��x��}��(y�T	.���T�͞��h��X%�=��=�I��o�3+����r��l+�V��WZ��=�d	�	���5����������2̦jF���'��r�_UUmZ���k!�*{��]��%_�̕���������̷�g���[u�/g�/�P8Rw�[��!�����u�|/���]6��ê��ǀn��q���5��E��tK��ǒu~mr_�+Ⱡ&WT��$:z�{�s~C�ו1
����ϗ�����c�E�c��
gŬW�O�Nsu������$I˃ϳ]�l�tk.H���7�<�}�x��ޣK&R��-�JY�[cH;�����r06�-OAO����3�O�n�c����?^yQV)&�`�%g�B�U�[FP�5Y��|���J�� Q���F@���P��v������|�6|�b}~պ���S�2���/L�ɡfɃ/ �+q��B��{r̆��{`Sd"�/�Do���c�y��XnA<�����CJԎ��3���P�L��Mq�����ڬ�ZUO�q��`a\�A��)*^��6mJɰ�h�?vVk�%�h�<�4�U�幹j�<�k��+q��\S�7�Zh:�0�#P��r��w�@�l���c�)�"}dEO}��-�˳&�R������Y�����>�LR(��t>��;�HyB#�@��������'�1 �*T1�MC	�q[�ݍ��/E~UE�z�o:���fw��G������)��K��)�D��IM��۩��D�1���Ӧ���}�%�5���XG�k)\0Jw~���,c^S�= ��¤���ڨ�>�3���i��8<��G;�8W9����g3��H �FXN�z�ݫjXt`߷���z��_M�aoi�v���m@db� H��H'&͔��(%
ƋonKBo���˾+�

c����]� &�¼��,_��1�Q�~d��A�Џn�l;�������>P�ᶕ#��$9@��mOH�H��C���c3ۥ�%�
A�: �������$CS�[f���0#v
J�_�V�
��e(��1ڛ%��$Q�,�A-�V~��^e�}I����7`�r�/L� �{(��N;�[���Ro�%޾oQ)f3L��k��a䓦s��,N����	��a�����ީ����Ȍ��A��'��-�_!(
%���Ķ���y��i��A �8{hX��n �3����c�wC/U"�p�	��C����>�����H.�>5���yL�>R��P���t��=�%v�5v��������7;+�}V�M�F�$e�n�*%F�F��ƻ ���$�!�5W���U�����P�6pˋXx��5GF��r�V��n�-t��یƕ�+�s��h��T�9�V�tAp��@폇�=Ϫ�.�3��R{k��Ɗ~���{z"�����T�T����R-��rnUG�H�v���!��i7����8F��4x�SoPڔW��h��*�bNc�_1�J�m�!)[vد���Y.鮰�z"T��։��a*%�X|�oZli\���7�ӷx��Xt��i�� �zm�ޠ��(mY����5>W�3qbw+�}�V��/!1T�p`�9�$�[�4"m��β���O}���P��%o ��Ϋ��sV��Q�q��fx��2�-��Wl�>e�˽�rY��f�6���\�d���yY-B��XvW���7��pH$
MZ����B_�",����6qVcW�)�}{�o�]$@)JOJ7!5G;�7bl����-�ډ���aѽh��1fX4q ��IO�W	0����bX:2����։E�r��$C�m%�od�d	��ș�F�E�^�d���bJ��i��vX�*�����	C��2^/�K�G��{�9�o4����0�v�B�*�E1��oJ#�٤~��.�&��mw��s�W�Lm��kʕ|k�W�^�ˮ�A����b'��Q�1L���/n��9r.����:��`Ef�eE��C�n�?[���s�#T-�C�T,Jj�t�r<���5��J3�#�zw�ʏqW��>׎�a��)F��|h�����~��	���U��K|m_��z.~r��B����}u5�0`S�kISk�P�Xvr�UfW�u?JL�q��������6��z�qF1Q����p���s�gS��Շ�s�Lg��=��=�3�qF,6�?#J�h�g�[i���.>{nw��(_Nh	 ��j�q�l����>_�)��-�#څ��ÀHLA"<a�4�wȒ�=��F㈃h$7́%C:�A�ߧ�� eY�(h��V���C�>.1�'0G��ȸ�c'uSo��S�{�$����F�.�E��ھN��ԩx+.c�ƢJ��0��=�u�F��������`����9�(�� :ؒ�������=�����b��\���h�	���jb�(�l6�����S��g�Li'�@Ϧ��LD/���PAR�W��UT�0��㔕��*"gr��$��@p�&5��h_�c��D0=z�{1?u ���
�@p��JW��t�H-A�S~SA�I���؟����ƀ*�yG��A19��Q�دt�/9-�(-�V6Nʝ������DR�:oW;/�JE����!~H��y;���-��#����P��:��@/�������O�#9��u�0'6