XlxV64EB    194f     9c0%����~�n�D�*��\̆�����-+O�b���n,ڶ�%�r�Gye�����>�s���X��4�3(�����G������c�m�J_����2)2TH�B�ARM��*��&>z"�v��$���@H�-#_��کsX�J�[v;���;��d���k^�܇"�X׾A��K�-����(0{�����<r�Ӌ���̐���*�b�5�=�#�|�"� ���{l�:m�&!�e=F�|u]�e>�9Q�>���|�ۆ���£L1J���T� B)���}�)e5���nhX���A��li��䦋p����V�ȹ�)a�H%�0���m��(8��R��\�jL�v7O��X��������*��H����]����*)��P�{��eg�;���>=����f��N,�xe��ndtiNɐ������<�?��;lqys3G�<�Ne�f���{��2������$��d�]"k�n��aѣ(���)�O9�Z��DY��s�8 *�86�)�7r��;�h@@?_�-�:R�y��{�3Z' �ˊGC�W��M�D���:@!��8�9},+���$C�zm�Z[�(�^�|E�~���R�Wƅ �2`�⟻�Q����=���k�(�Ybd��J���џ7�2x)�#i�� z���~����HL�5���BR���nF6)Q�,[�A ǵD�����?`��L�(���
���(���.8�?4I&���U�uQ(0����=��0pگ6��&L9��c��o�wh�������$�Wt��>�Y4��I[�MX���Y���c��+N*����?�Z�5Z�q��Ź���o���h��;Z8O�8-�N;(�v� ��2��m�M�U����l>p���"q�_��$�f��{�=P-�����s��y���<Id��hW��m���PB��e���Ne	�큷Ӭ����Q�x�%H-��<�GZw��b8����k4�=�2�o�<(J��N£�l���'em�)'�>�=�UJ0C�	}]�i�SU02���c%%���t*= �π:�̪�JH��㧻ds�J�c��+S��?X���L�e*�Y��	�q�=�nb�U�S�����ȱ>�m��d�Z�lAm�0k|�����	�^��t��;	��T�XY�O���E���@��r��ҷ� $��!������A=��bֈ�+�s�<2����ii��{�$�$ܖ��&����BX(!
1����-@�*��uh;'e�W$8Щ��L�:%�iL�	�TuI��f�`��CPM����0�F��0,���V�J�|����1���Ե0vd��(�=�g�uܙ��}ɜ�B����DVIf������AK�mE�}�L���G�08^bn��0�L�.uM���u��
r�xk8^�AU���i��CP�����j^	�-�+o��'6j.��G�lh�������K���6I2�����$��b"�˥i.�m��\�,8 �a�����o�4j#����Gr�Z�%��jf9�D-��		z�bK�4#���K�/�/k������.�WP�D�Uo���(�6&�	=EI���h���T1����P�^W�M��v]�fX�CX�/= �Ȍ8���ϲ>J�ɦ��(-�w�N4��>:	RX�~z#^�8�Ly}�u&!��
h�:�NA�0���IX6��7W%�)Z�/�G����:g_m�z]ƃv�$W�����@D�&�߂?wQ��˴���l*���tZSq`})���E0�pg��c���AN��Kâ��T�ɹ���k�a	 ;��M*��&� >� ��&a��"��0b,�;[�o�"�	t��X��1��^���ņ ����`�l۩�e|�慪�V��$"H:��Cr��KYQ�p�ʓK�k},�2���퀋FԚ�����/)���|���J�mյ�|_�c��
ޝ6H�Vl�C��_���'��-�;����n	�N�����*���
Mo ���4h`��> #<�Di���GJy� "��@ByH��(��+}U?��]J�;f�l�3��vj�Uȫ*ob����M�A���ʗ��Q�;s���2�T�� ��G�p,�<cu�KH#�o2�+nr[( ��;˛�I�FI�r�\sƠ5nud��4 �u�o=�j�/o=Og�,nzK���'�B�+��P�/�S��4�9
�����̴��De�W =´Uk,۝��)z��J����7�p�s�m�/A��Hˤ�)��cs����{�YS^��J��ƌ���>&�<����e���rcz*ƛ�S�3��m^�m�ȯ#X�nͻp�5��h���}��e�Ӑ$�]r�\�ڀ����G���*�m��h�';���q�Ώ	HQb��~�ɻ��8�e�Tw��5̝A�
�<��MB��$@���ί��_l3����G�|�#�?��