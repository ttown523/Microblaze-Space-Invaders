XlxV64EB    b718    1be0��5�!}C$�ʨ��
�Ql��j�P�՜��l�a� 0z}��\_�D@��}�kZ�Z1Ş�Jn�H
siY�5��Z�U��_Ɲe 9VNt�J�+T�(��h	-""<�c���[]ZH����a�Uɇ�ǋKC��]��m��Rj<C������V+#�B�m-hy��0M)�?n*չY��e��XMMsl�N|t�d�@ڳ���c-�k��[b1pT�d ᙍQjN��hi��l�sS�u?hz4�+�S�j�IɧT%���_��};��&PB�&j��%�xX��܀I�2$}�|�عS`����|�`:���x��z�|�9�/�|ȟ�ȷ�m�*E�}�Uz��,��x�4��֪�ī�mb�t��o�=����x%[�U�⭨0�~L�i>
?��̝.%�nd�q�b�(~>h|?L��}�_��dt�ާ�s�S$�r]T��t���	_��P�h��N_����Wp!�[�}���Pٶ�v�ړk��b������j�tJ��4�<ۛi�U�s��6�Ţ���OhC�vZ0�R1kD2+7�C�b-S���y1���������Ҿ����9k3}�:�r��=~�7->!~�ؘ䎽�-��x�G���}:�ad�T�ٺk#$/M~w�O�l����:�I�I��s��(�%�|,�o�-��E���`�4�bM�X~� ����5|.��TUX���ƿ`���J���u)����i�tz���@^�=t�LH�1������xA�a�y�ߙl������V_4���oև��W b�̴�Z�z�3��Ԇ�9[��H��;»0�8&�A�G�*�g���%�^��K}S�`oA�Ld�SyFHQ�y�H�	��*!�9}�ӧ�gN|����%��aL�d�<�1 �-u��&@��6���z���&��}[J�}����o�Z���hI������e&aQp�vu�fI���/�إ�@����6�`�!�%P�Ҵ�7ׂ��ra� `Pu���]���=~���WJ� Hχ�˥q3����t ]�q��hǛI)Jh�E%s�:�L�c�K�F�!n� 5�o��ΰ9�5/�zJ"�+��ܬX6��G��B<���Ӭi���*d�96܆yr�n�{����I?7��δ�1��2�H�&|l]���oHǪbz�`؁n%4�K"#�qt��T�4����h[,�R��+hIG�*�79 ��V��b%~(9��K�tݵK������+D�9ޫ��ۋ	fDH�����~A4�c�w��i�)9=�ۇ�w˘���W�&<7c�~0Dr�u|H��� e�j�1b=�a��p�g�=��U�s��1�݌P�F�D�}{_'N��VCD+��:��]�n,��%����d~69��(3�f+�ͥS�ޘ�+��>5^�2 -=4a�Eԩ���)�j�Z��<��x��_�y����g[��*�>�4�9��I��r�A5��XǶ� d��Jf��s:���_d(bƣ[9rV�Ƅz�뫅�ۄ'��x|P�)�Ge��~���/�;�9�BLv
�xN�A6����[�� ��b�*�Z��}J�_�eWt�T�ao��p�Z�<��n`�����<���wxNM3�ӑ]��MKrp	�×]��d��\��;N/<�ԕ�n,쫵�h��.n� �������ɋ�FE9�W?!]�g˧
RC/�Uȉ��<��CVf�"Lg8ܝt�y��'��qd)����Ϧ��P��5H�'ƻ�@��U�w�C���0��x�����'��M~��뷇�>/�ɦ�������5ݓ�z�hbр@�C*������mOa���a���8J��� %��'Q���������˳a	{��Pۼ��:WXQ�tEN���e�{C����|P�(R��v�~�N3��|[Z@��2e< ��+/�c�I��^�B�H ��㟸�4��\>y��h�wr�����jVo�"�D1��0�3�M��#�l�IѪ�d�;��O�Un���-�h��a��^_\8B�nU�!�ter��C�,·��Kփ�]Qq2c\
����h�9�2W�"���um���l#P4p�֒�ƽh�z1Jv6GtR?4�٠޼��T��rJ�#�	�-ɻѓP�����N��(����(�Nփ������J)��T�U��0��f�|:l�ve����oT�om=O�Й����i2L�l�~
�2Zt��8{֫4��Gȡ�b�"�?r ��|`�[�<�.���M��V�{�x<��Ϡ,e]�	M�e���y}:O�G�C�oj�5��)��75ܗPZ;��b�o2V��GQ�i��n�24c�K�Ҭ���ȓ'bMZ�8^0Z~W�ve���k,�W�t��NFԼ�}�3����Ԭ2o)�(j ��X6��"hb��^ǫ�@,?���>���(���z���!��$1< �"xn��t��fc�H�ͭR,��+����# E)�om���˴竨�dn�G�E*Rq�}��<�#�=���a��.Y/�Kp��g���#�UC�ޕt#s�j��G�3�'�*Ʊ��V���CrŽ�R}|��D7���+���✶dEX��Omkq�*8�}ۆt0�gz�n�������F5z�TϦ��H�7n/4;ʏo�f�O�B_�B��/{��@�m)۠�M����Pj��K�c�m&zXn6��w;#s�LKhJ���H���-
�w{]�=8DЫ����U��&@t+2��ڃ���t�U?�{������2@(�ڑ�,��fv����$�D��x��鮻Í;O�U���آ��9�i��L�p'(��h�
��A	zދk}�is�Èc6���������՗,�0��Z@2�y�%&��OgWh��ъ
�<"f��˥�m��!m�8��Ԏ1����ɱ̼#�ҏ��}(2
T��>VqE�M�i���>�G��&����h8�n�z����|��7Ο'Wx�J�O\��C9���b��1���V��{�� W{��h,ޯ�J�����Bf�L��x�{qչd�}	StE5I6n�,�`؃���8��~�Tm��C
�l��B�//�����Kgke�-w�Ƅ�A�h�/�6D�~���{�!�#>b���ן0�'Y~ac����c�Byv�L��y��ei�Ѱ��11:�<�����(7�h��r)�c�M�SG�B}l��\�/5i�����@���fug{�F�ؚ-x��b��6"���9fY�����i�ϊb����܇����Xz�iu����d��g�(�[�5�T��sӀ
�Rx�U���,?}�\I��E\ �W��D �yNG.�刁�zi:��C���aӵy�8
)��G��4�>��4��B�{�̀z��r�7���/F�D�����UĽrly#/�{ւ�����57M�S)W���+��	��4*t���q	����4�F�|��%�6g �����T'�zY�R��YR��9s�N���O��|�/�\�-嫮��f��i����`Prf��Z�-w�8��Uoo�m̔
T!+$Z?���OU�<~�x���j`U��M��X�a�a�L�=�s�<C���B�r�<s{���Ҫ`���B�COr4�ٔ>jJ�Õ��K��hN�%.hW5ĝEG+f�͈�~;to�Y0ȴ1�������U��5N�v]�ŝU-�E�2�b�G&K�RU�^Z���duT �0��N���X*n�L�+$��ںl:,�e��� q?X�v5Aօ�)s�L��K�n���ޙ/7O{�8�)�7~�R��b��)�mD��E���թ����5��<#������Y��%�n���������`j�w(n���ST�F���JY�P��C���GzkS[V?��H���"+�=��O������D�=����C�u�z��-��ei<���J�e�C�d�G��Ea<E�q�<�e(
�"��+z�.A�l�x��N���J� ����"�Z��\�SC3Ŭ ��vm�X�@7���趠+<���II@A$ �y,%Q�;�������=�]l��>��b=F?l�H�����r�<���R�/�"ez�lL�U�&�j��TJ�ߤz@�Θ�Y,\������z�T�3�n��lh5S�פ|S������+`�rWdi� ���
X�Y�Ue�0	PTp�HRMf��O�c=o�mY��#(:����+vHT���Y�1�MhX]���k���ڇg-����,��j��_���n�� 2)`LT�4%?+y64�4,�aak���l�Ls��[}�^v?�_@�� �l���I-]��-�o�y[fx8�qd�![�J�S��c</Ռ�:S\���E���|���iǯ�bZ��~�v�M~�ᶷj�����$��Oa�8.�&Q�Sz܀Qd�s��v��t~�}}�����`��Z���SF�(��k��!�p����0V��1<ox�N1�G�^���]��hU�X1�j�/�nMv�#����i9}O<-�Qa��v�f'}��m$M�iH���sc� �����є��,Jf��d4�^����r#]G!��g!)Rφ�u�c������}���%�����}���ť�[Ԛ�n�$�[2��U�%����[I��m���ʏ)��W1 *�i)Ex�����j���� W�'�{�6�E�R�%�� FM�����1=�B�ʻ4k�~Q���4[�'�[k�P�tx�>e3����r�d�{��۲�Zэv�+h�;�(���4K!R��I��Yڼ�U�2�{Cmq&���tg�I~-X:a�G�&k��P;���~ÿn�� �L�s�7�Xǒݹ�ѭIU]����^j;��V�����-��i3�j�J���4G��O��v���^�� j2a��cX��GɃ�u��ߙsƥw�ւI�Gr��%�,�D����r]�1�AA�+��nC��\>'U=s�X��K�]��t�<c�\7L�ϓd�>K?x���,M�\ tM�֥QD��~���L<g< nbv�w�o����~�����7���_�EÔL��#�霫L7a
�-���x�d�xR��lJ=���}�Ff�tv�D��2��.R�f��"$�w���r��  ���:�����q�S��Z|�
���ת:�E��Ep�z�V�㴧sP�l@pb���^)y�#F���2����Ŋul}��s@r�%��(����CJICR;eUak��0��P#<��aَ��]�/e��������d		7� �����\86p_f�������]��j�dUq��.� `�[y��x�+��D�aX��3!
�FPB���q���qD>����rXa�s!tA���*�%�h�h[9�C �G{V����$�/� 2����B��\r���A`M��LMN��DV8cA��`��Ү��wB��w+�׉��`պx�#X�K�" �뮁O[E��H�,T����x/E��]�?^ndg�_4��'�$6T�7��&=���0�ٱ;���H4��
��E����-a����gD'�&�rn�ЄV�(2F��?�� �՟��-r�"?a���M�B�Ӭ��fFȚ^��H�u������XZ=l�8�A,�H�3���X?��zÑ�=5
�eF���d����̹���0�G��be�`pl*j(٭;��b׋�Ĕ^�}��Ww}��� ��.�p��r�χҞ~!�j_Рd�����U�;�(2E�fp�/��6"��c'��KD#��Q���喩��-B=��=<�~�pO�����b����ğ������@��O#��p4QG���6����l�}�#$l��/+ƹ�p%`��W���y���N�E�a�=��"�Rl��R��B�6�5����+�{�Ko�)w���ɓӺ7�}�5�G����>��"Ӣ��/��� !��/P<��l,rhy��'��Q�0 ����"?w��e��&�I�Xӄ�N2b��ݣX�
ԛbk�g�|�"5�_�m�ˌ�븘��ađ��;y<m����oW	1Ҕ&�9���,�*�8+Z�̂f��s	�����l̥�Һ�DAp�����M�z�S�!���3�{��5�n[�l����ƐQk�F�V�Oˏj��ꁩ�B��M��#���֘W���6��܅g�PJ(����3�&Wq{��J9A	������.swT���D�դ�5���^�ul�BJY�_/��:�9Q���/;����c��Cm�F��M��{a�����'=Y�e�	��|4�y����G��̛����w�1��S#��֦�����	Ԯ``����s�����4�X�޽4Eh�T��6h;�� ��j���.|�c��z6��q��Q)\���Kܸ�5`m�����\E&q��}Z�,�
l�0LJ��n�Ƨ`�����+�Q�1;�@Yr�^|����~����j�\� ��E�E�*鎅m�al���H�8����;C��=X�DBv��
p��Pz��F��7���K���r�_�f}�T���D����f:��)�9Α��I��[�N��aRgT�g�V�`h�@��c¶)�`[t��Hqw;R�Mo
<�-m�G�
s*EY;!ƻ��[�-��{H+R�����b:ە��i��k���p��1J��ڑ�*��R?�}
�*b�7�m^T��Lk����e�'ݤ�)s�(y'��THjl���t]��]r�!�FK��Ü�\��<�_3h�~�WV������1E99�k�l�S 4�V��XkQM
A�p�(���ӂO�(3��_�0���B�����ƀ�6l]���ĭ��p���fW��句�*�Lț�,�>:��ޔ9(�M`/[��j�fb&_������u[P'g7k�7ښ�YO�wf>:�k4�NL�j��?o.;��s:#a'��"�f"T~?�%���1J#CH'"!��@?D(��1�=W�@�^�ËNba������5�����Q�M�h��*��K���D_�B6-��
A���(��-��-��(ⲣ��*B��:��>ܜm_�O*?d�,g�x:���W�