XlxV64EB    59d3    1410��j�W/5�a܄U㣉"ا��='s&�E�
`�j�����t�,�+����U�mld�Rm'�l�SѠ^Hl0WN ���-!;�A�z�Nt�w�g�S{�g��7���K�C�o��&�����6$�� 76;�n.�%���xBa{o�y�܇�
Qa���v^�,rO�(
�\M�uj �O����
C4%d9"�s�L];���J���)`�~Q5=��|N��!�2�q���\����Z�7�9��k��g�*��v8M^Wl�=�����d�=E��|�1��I4"�>�i@���D]E�7��ri(��~&!���%�{��u�K�����6-W!͒ ���@XHA z�Wg�-(��1)q��TvY�R�:�� �=:�1�"٫Q����:����d*T�d	��D��^�(}�/��'�^��Ֆm|�"���w#۫�A�5݇�U���y�^�\C�*G�y���`��$�9����{�i��?lN#|E�<��m߷O'j��������c�]n�"��'��Fbu6g�$e�z[��%�B�,����y�5*�	��ܾC��>�ʏ�=SNU��?�LuS����������~k`���hJA}	��)����.���ϰj��v�K�=m�v3��V��؁�S&v;�����3_u��"��O�r��uL����!6L<�o��=��C����!�p
l�&��x�V�x�Q�����Zvs���X�Ϧ��;.��v�1�/�d	�~�JA[ػ"�-���)D6�졋�T�n�BV>��xY-����g�{2|����s�L�1o9���G������7O�P��;!���K��Ϲ>���>��I젅���U[?�0�T�,+|!:|��q���^.5�s��q��|p5R�v��p���C��K��HQ�jB����CE��q����3��`2�^��3�x�~O�4��2R�H�"_���'��J� 5;G��a�t���d}%I_ S <���g����o�A�1�E����"�V�ti�MfI�T?��-�����p�|�r��z#��%��0�T��;>����/�g��AB�� �w��e
��M��Tۻ������C|}o�y��B��Y�3�PX&)ۨ�)(�:�X�9|��90_2�&w(�y.����wA���^���m�YS��F=22�W�����iA��p�>���k�����F��P��s#5�(�Q�{'�Ί�p1#M�Bn!>��I��_�n*p���������x���1��M�?V�I1\43��.��:%7�e��X.'aΈ��:��\�>j�kC�嵺�4ȶ!��ﾉ"��N�������-Q:�wOt*l<�����������m<��%�aUs�m_ժ)�?d�l�G��!c�S��)�K��G��?P�o����ifd_�S�
�U�bb���r�5h���u�s�Doي�I M&\�R#.�!ɢ�#؁���q�
�Sa�Wܱ����o�w�v�F	N�gheYGc�U�4}*�"��e@ȥ�M^��%OO�@1e���}F��z�mֈ�N>U���v�^u�M�U�p�ל�	H�+�^ ��y�:�}��0���p!BY��T����h����Q�2�\�ąG~��b"@_���[̿�/g�5]Hb�:���u���h�{I�'"w��I� q{0�a[=X�	�l�[�KVs�Jy�����*h$!a[;Y�-ĕj�^A�펫5���RD���Ho�\��Y���7h�V�������l�2$���
u���
ꛆ:4�0Ѹ*|�S)}=�r��S5T�W��,��~FЩ��/f��P��c{���1X���R=B������W�R*�3ub��M�6�qE#e�h%\��2]'8m��"6���K�7�Q.��Z�~=[Q��[k%�DHMTa�و$cY��]fY�¡��(uz}B�6��:�������XBp>n�+��\��0
��6��5BM��sh�7�$5���9%:�;�n)"�O�X�S�<�<��#��nta����}!
;9�B�Dl������]Ė����mS��mQ�z��Ɏ���g�#�J�b����k5�4u�(�K���Gn�CR��>D6���7lj"[��a��\V�Ǭ���[B�,�4"o���%�Y�zTg�H�u��p4�q� ��.��2���Pk䰲��ؖ�)(��'dw_���jM{��;�n.���B����]���6�I(p������W>Y��X�L`��H�������@��08Qbك�U{$�B'�C�6�aJ�R,Ⴀ?�k����L�C���B���������J���D���P���0#g(s*;i��;	�c��<˕�t��Z"z�]F��0��Ila�� ٟ%�]y���JK�Ul�KB������Qo��א+��${*����a)��ʆ����z���)��1�EYy���$9���1�� M_B�+P�aBiC����2@D�7��An��T8�j��s�r���}���T	��&8��&�ޖ�
[����\��p�"��{�'���5c��e�~�Z䃏E�E�4*;��FaH������θ��$�LDmٚ�"��Q)8�b��o%��{����î4�Ft*�i�.#@��' ,�G&���9��~Z��V��08ʓ;!���*�������6?5���R]��	8D�������*A$�̲>��3"���E]ʚ���k?�>x����<l�֟��S�Ϫ�5Ҵ�y����s�H �cҼR&r�jq;�\CZ�أT$�]���9��.
b ц���Y�7�i�[���Gd���t��g�e)z+�̳�i;�v|�5���<Z�e�>�Ax�Q�ɯ}B�d����g*J?OBK.5��o$8�ő!Ļ��1�Q�(�^+�[������[���"RR&^d+�F~�To�2Bj�_E�	)=�%���h�~��A�-X�}��o�6���熕��a�2g�SQ���y�5��zu�˪lN'�8�?��X���ʎzj`�X�a4�.0Uj1��iW�d�<5ƌ�L���@)�[�ZF��n$r��q�$�0,�=k.��wvK>#�t�V=����KVA\�:ԍ��������m����%�
�Q:�n�'5�s��#F��4佤�S���S�Z�k��
R>�'AtN�>QZ��/��E�NUٌ��H��`C0�+[�����2����(�%�xȼ-�q�.�Q��� �����^%�*��b��G�������C�:E�L�'��̓�r��U�#���r6�w$(�ý�N�yP�Z� � &��|�rV02vTh�u�2y������F���R�y%��S�.���k�e�-�{/"=j��yBJ|��[<Q��|j�{�����.�za��*_�>о�u�='ͣ���$��Vԝ"�ҹ���1+V��7ٚlXeQd櫄���d�z�6c��s���L�vbX�t^�d�0Sh�$��m�Vd�P�Lξ3xw]��
������÷	��T7�JZ&�e|-$.�C]���Q�m q�������%�"q�f�H�@�	|���Ǖ �p�҆ƍ����)��pL����M��^�>����tZs��ڃc�wu��L�V��e2����~��ӎ���r�PX%=�����`=fH�H�s����ƑiF0*v�<�[�{������r�Bs:C���
FPT�"/Z���-A3�̽��Ԍ`~H�b��k =�i��G�{�f:h.z	�Q.�L�\pr
8��Sk�����f�y,-��a�c2���O��w�+����ު��g<Ut�k�!�-����[%R�(S����]�{i�?��ڈ�捕�#��r� F_���)�	Od��:/�;�E`�-R~܏�qp�(FZ�V�'��9�6�vk6bat��oe�́h�'ǩ؛�Ƨw�6��)*���7M��'3���"c�um-n{n�c�.����)�A��e��AC�{����R����SÎ�E�g�	Y)�ʋ,=��d���f�͛�S �\��M�T�8Q��К3���a�5|� ��j��ʌ2�(�$�5ɦ�������ТA�������X��D8//�'!�ZO�~��e��U���cG�l|>��6�M��l�|����k��RG�*Ak��y8.��Y%�ҧyaaa�~�L �A��L�w�`˾m�\h�=����=���.������iixm� ��s�:b*$����)+���/�%#��閽��-�TY43ܣ`v �������C��-H��i<�d{?����I�W����jV�]�׍��9UtJ+��B�����W�?����%�nk:}�pYU2����A����+jV��"V=��Ksd�qVl�ƅ�3"z�V���&�ڄ_�g�n��B��Q�R?�hp��}����u�4�uVC]er&���HeTt����^�P����H���ؾ~�2�ј�EG;q�I8q���ް=,>��	�:�yK�CZ>vw�B$��%ŀ�w�;db>�_	s+��C1��Qf0!���7z��͚h�Lz����� �.b���"�G��{N5iH����AT�;q(��eq�̳C���}�����X�Fб�X�%�p�DeW-4�w�4�#�h�/sK��[��-��̇VZ'jTl��_OZ�3Rʀp#%&�Z��d�S�d,f��_���,&�����?�W��t��N�oյ�`��{4b�rP�bm8�"��՗u���-Uж�ȴ���y����F�I�.���SN��9��EU66A���(��ϱ�|!�Tv�����FRs��$��YD��svj�������$t�K��s �Ϝ������Ź?�ǮGFtؚ����3�a8��T�ӯQ�2'���e0ϭ��G
(�\���M ��7��9���ə̤cʁp#��6���j�/�v ��z�0��ǔIkIm�Jj�mh��~ß!\J��S��l��wыW����!���TۼT��+m_��������4�cf5�a�0��jM挵~4F-Yc��e�Y�)_�