XlxV64EB    24b5     c60UJ�?_��X�Գg&J<k{�k���;��+e�p���6'5e1��)�!�7���L�7@��W�}�����-9"�=y�뻬翭���B95)G���+���݉�է+���jη�~uo�ny�2|0ߔçˁ�$�E�/;��bꊔf���N��}�R�A>Ҋ&�Y)������J��+	DCx�Vn��zܻ��A�ؖ�<E�=Kn�t	d2G�/��P����C�W*�:�/�	[��X����N4���V�0j<G�P�s#�l����V��x��"7����[���d̳f��D�o��nRl��u��O��[��y+�R�g7����\�bEǷ{^#��b~���erc��_ԣI��箧��A����=�q����.J gA �F���$�z��g����1�:*���u'��b�Yi�AN}&6ò��GO���#p4��2�v�S�F�ٕg�K�S��!���5�L�a������������ŉ�e-��'�ܕ���c��LG9�g	���E��=%m�W�������q�R�s S|��*�8�K�fn�I����V��K£\��{���υy�]尛s:��!�L��{�jQ�~��0P��l�w~xa)�B�6L0TF�w L��b�5��UZZG��/Ty�4�!>��1�L�þ >0�X]�р('L̥�����B�ԩ�B�u�v\�$�N#N��O�;h{:x��M�r?@�L�TG�!�mٱ��j�����=ĵ�{�4u��vἳ��!fС�.��O%vEG|r7#�1�O�؞�
��w�n��`�kL^~w������g����i�<�} [�V�{�)y�-c�rBzg~��j��o|��e�<�&�)F{�(p�� ��=�-��n�9�7Q��s�������X��5
�ԭԤ2�(0���Y�6?9n'�5�i��Do�����&ϱ�,�U�]�K��Q}����Υ�r��Yi|Y���4�r�/�"�X�t�M7ǅ��%�ݘ�MeD�N�Iu����ﰢ{��U�&�I9��.���6*(�n��N����(��s췮�R�]��Y:�?����A\ɫ�,��95�,��j�l��O��3�)2����k�X�U���Ȗ�jF����<]s��7bT��?�]�]��v։���#�]P�h���L�����6$�Mu;��6Cx��g�Ɉ�Y���'���p�v�n�ds���ME;���"C,ׅ��9"��i=�9?&�\9��>%-�7i�YO��KaK�(��')�]������Bm���!�hk	��;�ᷨQ�L���8�z�5�;*��%�𿤸<:ԧ�+��irʸ+Q���eT�<2P�"�|}�ag>����.{��ge!Nw�͛1����7�����0��,�I�TxL�W�n�MA  ��_۰t�ʅ
�L_oŘh��z?ՒA�Ӥ['���(�}�됙m��d�"傮���&H<G� b��ZGP`�m�8"ƚ^���q%��fx��Ňg��yCм�Y������s�U>7Up�z�b4[?�i�Nx�S-������8ت9a�7�U9GN�c�e�����eح4���]�ex�"o���O���3�&�|��2��o5Yn���;�$�.��i9��lz��kpy�{�����$�+3��p{�I՟~}*���0e?��\:�\%��:��Asp���23W�oUe�]'��A�'����)mD��B���<��+�Ŷ� ZƦ�<e:��.����p�q0+�J��9(�o�a��o���s9�.R��OO�a'm�i��N��(=���k����� ��s�B_��J �A��"�ƉA�4bU�'���I��f�xN���W�����D6�X��0�W�?�t���ެ�2��mE��Ǹ��Ǡ�J��cg�z�'�|�6;�,�6�g�H/��kk�u���1�u@�Pn�r�ЀzZ8u>��,d�&뤴8�(W�n}�����U˝&Y�!E���\���h��
9��<�G��$~���$;�K�h繮�U�:|t�����#'J�w<�p����<t���-��y�ٗ��� �*R�"@����]Y���\���H�i��H���x��Jk�8�*�
e.tB��vW�t_.e1�-^��]F�F���a�)hR]v��\�`���u�]���8Cn_�q�����{8��B���|a��,!����H�� b�-�i޶j�@r\Q)TN�O0Pz����^zz^X�����PU{][�A��H��������J��~����$�ʶ	����t��K���Q���e�V����c�Bߏl�r�}��(r+���v�ڎ��9wc�,^.Q��Ҟ�}a\��K5�Mh\2������i�_�B~E�ai�FَZ�'�^�=��543oҒ�^p/�u+���/�6U<�DD{�u���ţ7��>��N�o1��||m6f�R�/���0JgÀd�aF��2B�X�}�YH�Rvg�*R5���Ⱦ�;�ئ��h�ݪ�?fFw�_b��P����M��8�'k��g�e�A�k&���km�u��~�^�K�9�J�0��,��"�A�n�!ϧ'trpӘ��ao����1���Y�����3�H}�n��J��ǃ�k(:D$F�/�۞'�E��i��Ԉ@��ŎA!tt˂��F�N)��2tV����Ǖ�u��@L�׋��u�1�-�S-)���7��Cv�>�3	���W�lQ ��H��4#3y�bN�#TAU7����ih�H�#��}9P�)�ojT���[�8���q7�i�{Q=��s
WVr��
.��6o�8��TY�]�`�h=)���O�j�2�{��k����7T����H;����"m s�w����l��$SG��+ Њ���A&Ǥ~:Ӊ�("��ƾ��YD%�U��oH�'%:��Y%�V_ɢ�N��!����f?(�/J^�~5j��A�&�R�����_�o��ϕ��ͦ�5gM�Ci��,M)���c�{�5��![��o6K��4�p���~����^�Q��ܤ>�"ٹ7����:����4��c��{�Z�%1%�ֲ	]���Y�;�i��/�2#v�NH"�51t���~�����,i��T'��XDi