XlxV64EB    576c    1410��O��}�
q;���Z�����Q�V���ڞg��SQ�?h�+����=�3�ѩL�����xO���U��m�����i(��ްt�f1}%f�!��Ŭ�0���,�M@3�ߢ�ϛ�Ͷ��й��6�^�Il$ɬ2�����2�Y�83T!��ĊR���d9�����OV�K�	Y"rHM�F�|���os�#�k�S�뗾��ח)  ="ϠR4�=�sC[�=���1ޡ\�]�?����g}�@.�je�@�R�e�-�&�pc��?yŦ$a��,���dt��~Iޔ�[.X+�aa*&��1"��.�V�K�J^5{kן�洳� �T�v�U��2=+�8�]
f~�Et_�\e-���W���!������e�X��!y\X�5m�Y���5qֽ�`�<G�2N��(6*,��t��.�5�u��ds9A��/𧋝�`�Ȕ==tL�K/����Ub?�-g����I���|@���+-^+�_�f;q��%J1��E������'���T!��6M��~un6����9���u�-�J5��\֔`cGQ�9$�J�.�*�i�	kr�&�mr�ch&�X0t"Š߾*C"Q���aוyd���%��ԢP���:�	HFtݣ®�52�f�ԝ�\aw1����M�����x�j��г����"�1b�=����C,�]}�6NNڅ�rBL�EF�yV��g���1��ZO�w�vql�88�>��j�G��Ȓ��Fv�5���tBy+75���\���)D�80�ݏD�pG�=�)��q��͋W�\~�����jeS�`v�S�6:_qo�<�T��Z��gh�!�+Ni�P�c�$3�1$�s�nH�~�_I3��җ�0�Z��7Vs2���P�G�DF&"��QG�sd����&�������L��������g#���XY͎�q�x�e�u�/�5�>v��;:
m��Yg�/�
����\�N/�/:r��'�{T�P��Ӹ�T�ˆ4cj��N���N3��ͫI������<,�^�N�g1l(DX�+)�2����
/�>4H|{�`�����uB�H%U Lw/�g�4�e�l�U��
(M#q���>�#��9�Q9�{�}���
���ɕ�U#�����0.�.�����fBF/��� ����HMKp��)e+ �D���vd��4�;QYl��VEN�| �}ɾ��F��쎇G3�'O�d��qN\�l�l��x�:�N89-��_oj}��]�d�z�ᫀx��8Mq�i�2��2�2E97�mV�􈱫�&B/8#�c�� +:��}�ܶ+��YA�_���XhjG6��0ݛ��Rx�Vi۵.L|�҉T��Fg\5D�3�6��Fy@�{ί��P���po����8��Hڑj9�xu�?�yU�� ��f-T;�X�?`�������\@����_��M��l��euH=�4Q.�8�v��Z�{� )�B5��~cܿ��\�j�g�,W��
���e�Áe4��z,|I��X�%-�����@k�	�O��.�H�ɷm����sCM� =�g�u��2����'��\;+� (]P)��5�mxNp(��\�e+z�Ny@9P�N�j��qn�l�6���M�J{az�6�����d�U��l����C9no$�Y
2K#�ւ�|w,Y� �:4j��� �Q������5���H�6�y5jꯜ���Q7y�����ذ�r�\(t|�t䤮0;���3�C����iza�#p���+6j�Y8�{�b��qp�_�w6���,�s!f���ß���Q\��i2o��ƃ�K�o�q�p� ,<'�IV~U�_��7���JD����.��6�����t�P)}6����tc��o��Ϟ�͈
��t�+�(������P��~?$w����|�VBm<jp*t���E̴�e(�,�"�����p���SH(#g��"cܧ.A�iڱ#�I�KtR�����f�*cjrb�C?��E��wj��y�����9YMFO{�+�0�(4Ms�	*��n�?
��!5�i�6� �pZ=�H��>Br�3�2��WS��R}�Q�t9�������?���ަ��a�$��#3΅�K����2=wd:ԇ�_�H4��%K�JGw��9���lv���"R��gYh���(�'�u�QL9G�[#����	���I`"s�C���WW�G�cH�����	��>ˢ���O�v�a]���=`߼Gt�Wl�����3��i��*m�3A�z�-\�/�U���ҍ�������#-�m�X�*fH	lj�=�e�Ŝ�cY�($�Lƙ�1���B?`�rcN���<]:V��`��_�|��q�+|oÇUl۰�(b��>O@�"Hռ�M�ys�K_#I~G����6��$��E����Ԉ�>{,�P�_�J`d6���䇩 H��eL��90:5y����ᦥ��iW(I5Zs鱇C��_�_�2�b������/�Ў:ק�4X�uG�_ɕ�r����vg�O�(�4�nXa�w���!���c�r�i�ڷ�����Ӵ�.#��V�v�Dz�����t�+�R{놤��n,5Y�ZR��mqu��H�D7+H �㟶�
	��_r�zØ��-��Z3?����a�-�n>;�H����z3r�ٙ^�EFu���Y@9�ӥ��Zt��߂m�%Sש�k�t�Q��?����	#˩���g���3��`;�f��yW��j\�ۗ&�6�J��SCnY��O��}�p����Ƌ�<g���OJ���-wv�[��}m�����:V�`Dj.n��&m\u���=���o�T�i0HO|��ML`w���<��/�r�	ٔ����3�]ԴH��0�<�����ܑ����
�vt��g�E8�c+RҢ�<�����.�P�M }ػ�,m�����PH/�U�V�
�fP@ݹ|r��
���U?�{�y���HT�Ϧ��`6���Mf�2�m�|Q�4�YN[:g�tI�L]1��6zɓ��� ������d@[�Ӷ1�Ǎ9	�@g)�-� m��f�L���-��e����,�P�0��n:N�:q�L��ь¿�Z>����馒SzW��z�&�9��-2��!��$3��[d��O}sѦq�mm�#����&�)R:�2��Ƿ٘7]�)9������@�?�=�n���f��u����K*�<%��p� @i�R���t�#-gw�yI��"�_��w��w
w�Ǒ�s�4�����E�>9��`�Y9�y!�5���$ok'��r�W���5�{�󵕛���$�B�x�ٯh:�& �1�5�@�-�㧆sTK`�woyE�P{�7�L��t�a1���C��A��V�����v�����9h،p~آ,b��4�v��|t��'���]�)d�y�*�xZ��Z���@���s1�N�lIoq{�ª�*1�14A22�~p�-�מ�����p�s����8!��4�|����?� �͚�z. D%�	�jS���\�I�SzϢ��M�� ðO����{����	��P�o[��������[��ۮ ��ހ ʦ���-�/ek�.}&?��[6`I�U4��4����qt��XLN$�ҡ�ڑb:��T6�j���'����];�<�K16��`�m4��T�5��Y�	m/��֪�y�'�!���Z�|�w��鵱����:U�ޘd�X����D��f$e�K����7aՋͰ���2����-X�.
2�<�h�_� X��	�ٕ��;�2(��H�-��
�3���/2�K�f�DX�x�_�����e���"+ڡ̳ c�����ـNK�5sӭ�Gb��5�������6PD��M?`��o�eq���/P)HPH ��p�+0�F�.�*�����w���h�.���A<�ziju3�=��gJ7��={�8������ �p^��Qd�f�7�ZL�J	3�l�k���s����a����Ä��^��	"�d���Й�>�m�y�����j6����b1{�%$ #�>�E�1O�D`ڏ�=�i���_|��P�~����7����[� �sC��ޯ	��\���RZ
��E�{m���}���z �x�qs��Sw�{uU�qaQp�j�K�_��F�}Ů����4��;@�r�ʘ����t����GlP��!�̱�ޣ:�~E�|F�6���!���7-�"�?��34J��=�3.�^ ���1f�*�Jq������җ�x��������@�HK�zK���'s�Kޖ����b������Zm|s�tv�e0�T1�Xi闢��V����;��2{J�	"O
/�3�tR
�{r?�#u����v����bQ��Q�^D�p3Nme�N�׵i��ԡ�m��J���e�G�_�Q؞ ��?o�}���7���׍k+З}Ĝ�+M�Y�>/%ix�a��°��^H^����;M����ҙUl��EL�.ϴ���8v�;��ꓡ콸���>�M.��}����؄M���c��:<���0g1�H��z � >$~=��6�eUQ#�<m�R	�ڷ�t�v�T��S^g�����v�[���+��p�) �5W�z�,��oPS��܍s�58�:��=�T��r�W�Ǫ$j_˅w(��C$�Y��$&e��$�x*�m�e�NQ��BD�܃Y��P�@��JВ�P�Z3}�ȅgRAh��Z	�����D�$q��!~�}�<�켿7����3������V��q�G�o���kXU��+tj�צ)�2���̹��>�V�uD2�������#z����Qǀ&MsU�~��n�x2h)��n�OʲlB���$�+/Ol�T�pdq�W�^̑
����x�Ơ)G��C�]'���X�C��UK3����[�E�!� ���<*D���P�5R��=٩�u�J`������O����phA܅�a�lֿܨm�"'-U�os�[T����0����e�%H�G�$-�d�A&���V�4�� OU
�_�{�u����{V3|�]ˆ�^��3R�