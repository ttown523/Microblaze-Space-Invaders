XlxV64EB    7526    17c0��V��=r>wޙ���a���T��i�����b���ק�"d��lr�̣�DŲi������Cw��*�n]J2�Nz���x�_"ђ����<�(������M�"�~xj�����=R�0	&�3�����Z
~mM��l?}�����rP)ʧ�d�~���i�.�y�;<�M�����IV'la=o#5;&v0��gOB�,�o��ybH@|�W���&�<�Ϣ�����7!g��Z�i��A3��2��Xn��.��;��������={xw����b�f��|��hF�4 ��}R�!�x/���8dP7�h����5�-�r<���yO~���w ���R�*��x,��&H�����.X�r21�D�ܩ��Wν������5;�0�`a�� $L�NUU�W�䇼9yu�~��X����@?�	�����-E~�t�(�f^�hې*u&��!(	��
0�
f����uP�����&��ᖱ��h��[�}��[-�ǉ��!^.�N��j��>�w����;!���o�R�zu9ڑXj��g��DB��Q����
�mxQ��_]IVȽ����{^�uܫ�����@ŗ>�p���3�_�� ����	�.ā�bO9�H*#5�jY�w�,w.�kr`A�^FC���൦���R��O��p�@�2�7������N�?��H�(8�z���qO��a�u�]M�n�{�#�sI���9Rx��s���'�Ҩ��j��r��7~�/��gw�q$~?�h��p��u�wD�;߮�h����'�%~�+��o�I4��V��1oC��٬�ϓW����D�,�Rۨ��iDג㞩���
�$7fV�_������O�7RY��h��@<��;�eJ1¡g�Z�߷�5spn�qRo�ŗb�y��i�JC����c�����:)�-�s�C�^�J6��h��@�&�x&-�o�U���|6yæ�	KB"��0��/t�W�:������;�*'C��d�S�G��� J~֤���'"�A��G�`б�RĿk��.�5���+�.$KZͼ� �utգ����U>>g�hCH�^�j��ĵA�M�I1�����y�?$�.�0�ؽVg|zi��i��,���U3�'�*�^�S�_�L�~bIϜ���+G�1s��C$���5T3�\^Գt�?�M��u��� ��#�i��,�9�j�s���im��@��#���[|p���~��]�y�o��P��
��'y!d=�B
��������@ݏ#dK�tR,�����}mT��%+c(H���i�+��'��W��ꉠ���+m��`
2��$�1��kJ�?���2�
In1���� ����T)��.�7ʼ��������0� ��ܟǑO��a�K�s�dЫr�=��gZN�dD+��	E�g�8C���)��Ș+���秓���X�X�D2"�#�F�AIȑ�F�jj��})���<]�)S�_`uoF�=F�a �Ky���|�q._ko�SI�	����+�}j*yߏ�������U�)^%��+��
���{��ʳ{W�1'����e��� �?��F�6�`"����|)�z���|w% ��=�>o��_!049.�P8.NB1��]��mw����|�\qb�3���������j�g=��-�ï]y0��*��nwc:��x�6��%Pd$���k�	M�bix��l!?Zr�Xz�'4� �.T�&�E:��w��}H�)����c�Et3�Ơ* ��Ϥ�|��0�'މ�ʚp�S�l������q�}����m�'�tюk��Cc%�`��Yi��
o�?�f��-������+P�c����N���.��C��(�oC'q9�&��h�^�S��a�MnY�� �06B�Xd�����v}8�U��[p9幫,%��W�3RP��D=��DO+*u㌨�z�й�6(��K�!YS��%S�\+��\$�3�B��[`Y�et7q"f��+eڂ\��?���A,�����R扉�A�t�#��j&��t�6���re������v��X�:U�E����'k�;��+��
�
�y�M��!�֓m��6B�jY ��l��������3:��ss�dH J"���v���_�^��x��[ 7ؓ<��o`M,X�g�s 0\��mQ#OXH���8:�0;��"�{��Y�
>�c�1�F��G�*6G&������ dYI����?�F�Ʈ*|=)h��g���y�rA�	�#:�/��
P^�4&�X�*E�%ܚ������$�Em�%%f �_q�܊���w��\Ϊj��찪:[�o�XG�5̅"���i��ةnV�w^U|:�/Y���#:�ȟ"@�iE�e[˛���?�t$#���<���[{�#]��!u��E�(�b�G$�{J!9)�Eb)�"(�O�����L����y�ۛ�@΋�t��]0�͓�#&}��@D�t�6�	Q���������Sf"J�E���7.�K����Tq�� FT�l%�l�6�vh�昩���s�Y��t�K���<&��<j�@?��s���TEq��"�m�>�>'���Y��%�#�ѰL]x��x�g�Kʃ�2�ҩ�#�x��>^�
��ک���6d��΄(=q����=,���j_c#Z� �J:���7���(r���&=F�I���o��@D�K������x�]m�}�_�/{�����X�w��V��z�g8�,Q'�̘�F3�ʕ���^��K-p�X���TP�%CS�<�r��(Uӄ�(�w�en�w�LF���*m���s?��`��\<�2�)v�w�k
��y�yD��c����!|�ׇ�����sO)$�W�����RV��Ǧb�$\� ��n�sjW�V�C���$0��TX%��N�`�lk�m
Z8p��GG�Ӆ|��������.i����t�1nM-���~U�8>͝�u�|�t���TV&��hX�c��'
 jk�S��U泮G�d���ٳ�U]j�\�7!c	[v�b��/1� �ݐ������o����z���/�C�0�9�{]��7}��"��q-��1�c���Zv���q�wv�G��d.u��y�,zY�na=u�0�8$�0*�O��㋗OWJJ_��q&Gz�?���h������X	�=��&U�3�)�JSG����rV����ҷ1��h� N�j��ʠ�:��8�v�c��.�[<Di���#��T$�WV))ە���)�2��T�P��H���\���x�J�{�52Wǲ���ƦE 9�$��rwGb�:��!���I�l0�H�ܦ�%�;+����?���O���ک�E��J]����4��Ox��D$W�T��u8��ͣު��{DVY��H��:e���Ļ��y��.�ܷ0j����P���b�gv��NnO/R�L[���V(�8mM�����L��|�.>HJ� Ĉ#�yXj,���+����D�<x<l���v�t���7���j����<���g�D��'(���3����wbKE��S[�ay��'�k��}���E�)ϥ�̀�i�b�m{�ZJq٘��� Sw�mE��V+��9F� �j��2��Jj�q��_l��?d'����)��_�	z�H�v��+5��V+���?�bTS�vvr	���"Kݝ��*J �A߱�����'XFS��&�1�Q+�`S;���/պu!l{��`q&�e~�,-)����vP���r�Q�:�������D�pz�]� ���͌��v�wq�y&�m'�s,醦`r�����N�mf�;���4����C�Ut����7���ث#��7�1O��SY�l&b��j�M����~��dT�>n3$���M6f���]�R�'���d�|���4o^�񝷊� uf���6z�����Ϥ�B�aU�g����.�k�2��a�$[�sP@�n��ϊ��G�*Z�D��k�N�ᶻ&Ĳ8�ٌ�r(��9�����㼲2�ۇj�
I�]6���Z�k�~D���fZ9�?srof�^��������p�]�������D'�0���)�Qvދ���6 ���f�ݟ�%5�'Vo4��)�4f��} ��k�wuy�P�/2w1O%��[̡n�6�G�j���v�����]��^� �%�z��|����Ԃ~T�Eo��ھ��Rj��Z��?c������ئ�T´$�4����Z��>3O$��|�o���	�+��n0�AIg�c���l⛪�d
�u��\�<����w���.氒�=#>t"��1�O�~�����-Z�����-��4�w��T�=:(�����T#�+{+۶�o�tTg�3GVK-�ޡW|6@��|��-��s�h�����ݒ!q��_���Z��y^P�n���rG�k��l����%�o,��&Ty�)Tg=��] �����) �Cg��;QY�FK�������N��^5�|$C4I�!;��k��X�D؂Ta��9���>E>��6;�qڻ���.nrx��VZ]�k�6��5�ᗺf:?�*~��+c_k16� �<U����g���u���ґd�Kg�w��Bj�`W�&B��?X��������)a6c�H�f��7�}=�&I���$��!+-w��@+k�.beG x��}���5c�_���w��#<I��R���tBn� Lv4�`MB�}ѭ�#B{��m�t��99pYq�GI���W���ȯ�a#!q�!��롩��=Bi��Z�r0�}UE	s'-�9��ч:Y,�r����~�y���a"�l���NW<��O��%c4mt�[�"���၂����t7�'��v`�1�A:�ӷ�.m��Ѡ���/��VȒ��.*�z ���gҀ: o�6[�2NhTMՙ�Ha�cVӗ�u0+�
�Q`�����u�2~>���#�o�2}+CNKiQťD��Un��w'b�t'�����`=M��"���C��P��|��_0�Fڱ�������8/��ڏK�[���2�6�OS�S��?��ɒ��sѡW¹�	�3�P���#�mOÈ��wKQWO;[CPf�|�)����
�״��5�tp]��7v��rz���9q]��1�[a��� �%��2�8��Y��H�Y�ߓ"�w�v@nn�)��ٰz��e4�a�@ɗ� �z�y40�<���s�wU�� we6�gҨ�@�:�,��x�/���q!�&�>�U��X+eaFJ��.A�������J����÷|,C#�^����1 ��6�)�U�V��!YĶJ;���9��I�^{B�C�*�M߿](�����}��Lζa�b?x�ǓZFS$���7���-��C~�A�E�b��J(���Gz��-|���l��cŲ����^}:;�e�����$�~�<�
�+"�˅q�Y��;�^�����y����X��#��Jm�/�Sm>U5 �濇Hw
�F��k����m0�$�����|�����\ٯ���+`8>F��Kf���q�*��x7�θ>����Y �PA㔮���x{�ܴ�:j����k�z!�Cf�iש[��i͙�c=uXw��'x�t	���{�.}G��h�d([j=D�M�n���1r}x�� �L���?ꢜ.RYÁ4P/���za�����Fpb��Փe��u6�^�&`W=h��ڧ�T�׈H|N���� ��o�a��lq���n�MZ1wBل��#���U��-M%��J5���¼v.���y=j8�V��V��"=�j}�&4��ڮIU���u���ʴ��X������s���Q��I�₰�>��n�4{�*T�y��r�4ܬ8�i�|]�����:�1�B���%�p�k�\����~#��p�ѽyu%��2�O���#݌ѡtV��S��v�[�Ц��K�$���ܭ�C1��~+
�=R����,`=���
�̕g�*ꮿYkZȌ����X�'�ѱD�K��@��%3"� �����,_��cn3�rw�