XlxV64EB    1ada     9e0�'�O��c�����'lq.���	���`P[,��9$����e1��W�׆��=�� ���ݶ��d�Sj?�w��/Q���+aʒcj�,����l�~.8!��!�GA��$z
���P� ���� ���!�X4��)c
�E�~�%��^�D��=���]{"�e�Ȉh���ܱXyh0��b�h�mE�L�s5��dd�=��!�݌�2�1���g�<DW(�K����R��rÁ����ڥK�HI��;�ޒ�ۖD9���/U�N�/�6$\�OLկ��/�@�V��9���E��CKn��9�Y��A��6�=�v	�*���k���3�{�WzQ����0N��-v�s����96�[f5���O�MI�L>�u�@�"1 �Q	����E��g%L[)����y��q�U�cJPT�� �lIiu��(i5��y�j�K��q�����o]�ܧPXE Eb'�O��ϰlG�l�N���N��TfI��:!��`� <Q��#���WE��e�JH}��nG���H.�o(�cAF�6�~��^K㥗��K5��H��#z���@<�;����H�0��Y7��^�_:��vV�����D��|�lߢ�$�2��+Pv��ƽL��|��'ز�����n+�U�b,��7�+�zv� �J��2c�rۖV���	4�W��t0���k^�S��ɗ���H�8��d�Ug9��B��%DZ\��v�A6��ǌ��	�Q���F����WM�G���	9�8F�� �0���WP������]�K�`�I�|k��䎦҃�隣G�Ⱥ�$�ے��%ϧ*�V�<�	��v� �V��;��CW$��9���䢞�[�,O����N'��{^Ί۴���À7��e;�31��P��0��]�2R����h�2/U-��?�ԡS.�l���<(�|��M00�@�T�Yb�f�a+]L93�	�
^P��#�D���� Ӽ�ΆIm���~	na�c8i�ϭ�a5��4R�,�Ǚ���.g�b��dO~���y8ԫ8_L�N[�L��{`k�΋6���%~���z���+�X�+�%g@��u"���ߵ��<�զ�Js�-y��@9g��1H��:j����!�͉�C��{��#_M^8�Ƨ|M5��U'*�n������WbS�x�p�+��`gK�G�O|�~�>�`��C�AwQ�#��=C|�xv�0�xFu����+���a}��)�R�d1t�E�n�Z$�}����m)�JH܉�0�#�ò��4�IG"���CMB{�`@�S3$�9�b2�7�1}Q���˶�&�����abc�XO��$�-i}V[�����ŖΤ����헨�����҇	�g��� ���% :s���7_�[w&*����'ҁ鬍������tӐM�Q��1����G"�ZO��Qd)�ȉ2��I�(P��[���c(Q�L�U�J�q�V����\�9�� U�L��Y#r;��}�|3�H�J�h��O�2�!7��l=�Q��C�N�V�����/j�х��軷�EΎ`C�dd�u��g���	�����b��7����Y;�j��u�m^8�UBX%}���ʃ�,�[�U�A�ΥG���qU��ꈆ9��`W���Iք��#��I̕ޮkx��嬰�E�CC�r��.)����+$%��!�Mvj�4�$��lQ+�K	_ri��0z ����7@�l�����v�����Y4����h�D�(�m1D/�����WU�<�Mp�0rؒ��d'�P{'�ԯ+
V�!�<��v�"�V�/���u���������	��i���&$c���4�U�{@"R7�CJ��r�m4��n�2�	+�̒��ѕ!-��
c5}#�
U��Ӏz��#&��H��8�X�׿���$���[6</$������Vb��n%�s-�ē��ű9���oU؛|�V�0����R]Ef�Ak9���PԻ�1�m�%��6B�3V����Z�S�A��w���r�<�)�qЄ�MUz4��V$ﴖ/��B��v�%�� X	�ӜlN��z��bn"��|HO���}:� ,gO�#n3��&.��Ի��?[��FWE��z6��^NW'��2�E�tB<48Vv�e�ΙO��A���*A�5�A��Sߢ�!���uN�@^+3��
���,�ƺy��J��x;�]�R?�����8F,�B=V�e<�y��D����T�g �/| �Lo���H�1_�a���c��zm�m�H�cD�`�[>�� Л�?�>HZЅ�����9p�A�m'/<Ȳ�K��C�d�c[O�����[3�4.�n�T������C�Ek���bz���V��l:�O���q'��T���B�;�n��F@�ʁv�+lڂ|��p����!v�s�q]��6����My��R�L�Io|��C������h��n7��Y��d�0����U t`��y�0�9f�6�	���#y�����*O�N\�ܙ��H�9�