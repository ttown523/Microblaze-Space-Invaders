XlxV64EB    fa00    2fc0��m�;F������Z�l,FIc�B��
p�)�P�o?ܦI�gQ^Qe�/�
-�L;��qI�؀�������A*�>����b���7Ɛ�����1�W�5ޅ��p�n]le��cl_�j��幮���r�Y��sK�n(�����dzlהk��R�EΓ۔���aE�ޥR
=0z�}2&�Тg[i	�4J�a���h�f�M|�[1W �A��|�R��Ϭ@��K��x'j�Fs�\�&h�����`:ck���-�w0[6T>�%�v���ǭG,�4Ux���<�M��g9�}�(P�`DB������1� �8 ӂ3u��,}�7��Ye-9��f�n�������}	�u���[��SNn��>gZd���6Y��e �P�T��,Q!k��ˀ3���r�o�]4�ۖ����\��d^�����y�jW"��C��K��6]$J�yB*0��'��K<��)�d�+"������`�3������lv�j��CMƂ�&�KeplT��t����f��x��\�3T��Z�W�k�=��F�.����}x�c-;�0;+� P�$E�꜡�m7%�b�|�c��t�����5ICT�I� ��{涒}��!Y�Nѧ~�Mg|�5�k��K���I��۰˹��/��˴ww��%�@��`���V �QZ���=| ��e��Da��H������iR�[�oWtS��4bT�Z1�J8h�fÍ�ӂ��w��C���l�p�T����+�/ݖCۇjs/7���=�D ������oN�iIϔ�'!��?�C���cK��1�n*�d��oDYf`�e���Ù���#����	����cXD	��gmܹؒڐ�N�f�K��vD%�փ{�-_�)��mZK����H��˱eG�K��:u�r�X�8��¬�4/Sn�$\�/
�YX���l)��;@��'*�T�MWé-O�VE�,�ܦ�5AKK�: ��:Ph�B��x�(�4J¸�������j4V01�L���֪��::@�'HT%��b-з��|.��I�v'�!_w�&��̻��!WW�y����6�v8]��g�:p�ֈ��MJgX
��̄B���i�
����ъ�j?��9`��ʲs&����֕�L�	��m,��ĭ�z����ȗhJhե�KĶ�b�jk���7�a��(�����A�G ���=�ey�.�o�݈�c���n]oC�R�K{/���/�1@h���v���b%]����o:��G#"�9pD��v��W������nUP�Z��W��2`�6�y��0�T�d����]9�0m2�����n�h�_Y���{%��<>)�/hة	꾥��3P:}zQ�O�k�d`Q#�i:�4��_���~i&��YU-��x��ܘ�K�W�8'�I��'�D"�?Qys_E��|W7i�����&�f�+��|@M���ȓ���aW�:�!X�L�dc=.>���^-hS���Y���W[���5{� q����z��u0r�����=H�����7�P)t'�Aa Gy��+?CT��w$L�S�H}4��Q�8p���洯G�@z[VTL�]��̙�8c���뇆�m�J[o��Д7�<�O��.s��ݟ���vR��VZ�_�q�}��꧓��q�@��W�c�{L�sΈ*�I| o��-	�na�ھ�~�l�-@�L8�r�!$Z!��5�'X�l�����7������^�����XϨ�DZ
����lr�pQ�b �8-�<聲�M�*�G�#� ��
�c�����J��$B7\,�4T���Γ��F6�ri��!�?-�)2��@Kc�r�ۺI%�NQ����K�qIӤ�?�q���D�ʃy$Dڔ��H>U����y��G���QM6��H�Q�k-̨�m`9|��1u)c�<҅D~0�0�3٭|�AB��_M�z�������TJ�!?S�a��As9\�T낳w]��F��B�>��v|���Yf���BE⣒} q �	~�b�����2 ��̳�Fd��a��Z<�?���y~I��e�X��Q�>���f��3�u��D�� k�e�{� '+�;��1v|f*nYO�;oW�Ϯ��pt�G#���<g���^?(��#˧eMv�8��i�H[�I�/�/��V~��h��a�gA�T@��7edRZ;F����9����+�u�{�:��P��\��ZSN���}��ݵ��f�v��)��j��g��̐,�ٍe�1�E8e.�vMTؚq������)�������E^���P�� ׏7�=�]f�����*^�M���96]�#4��C]��xS�E���
��h�����
�Z����<��f������I!�CQ9��{`����#3~Z��<[�QZ��G��of�і�ry��|jcE8�	U=D����(��:��Ƕ�p��cٻ�.�4t���^{큄�<�H��p����e�?g�G����	|��Ȳ�ak�g2��<�s�^n�7&w1��es4���UMota�f�s���Y�f��{�{Ɲݱ���N�oh�8B��j�j�:N�S����W��H�AP,ׄ����:@�;�g�D���
���o�!���'�;Q~�~.&N��
��T���e��Ut��+*�	�c�r��Z�߻�K@q8f��5eS1`�h�)�Iu���ͥ��moJ&Y�9J^��4��aA�b�kǈE>r��tg���aO�	�ZԲu-��0;Q�`R}�������Q��K�"����z �!��m���E��(pk�ɻ�dV��K(�-1ɻ��<��#�*�>~t%�ܧ����G�rb��-<��R�yp㈅�^��v���G�'g;3���)�n�u	����_@�с����%'7'q�՟��}���4�J��o�M녠{IL�5Eq�%FrWݖ�gp̱����� x4Ҁ'��y��3]-���\�EM�����H��.!�����%F�g����k�� 4�\M��#;�.�;�P�l�{�z��� �8��ڬ��$��eԩ�b���� 
����ɚ��V�Q���TZֵ��As>�yu��8�i}[H��Ӻ^]�É�O64u^�P�h��u�L��e���GR3�p�7���¨��Cf�J��k{�S�1c,�ez���4]��L^�y.R�̠�e7x#j�q�:�_J`�����nEu��\�xT�=���ͩ�F%�
�x��:�~DR�nyǤ��42��:�4���"�G�}1E�=z��fw��Wfé�5�� ���
v0����
���ØÒ=+m!4%n���C�p���a�KT�a5����w�s�Q��1��Ar�zl��wG�T�zϥ�����:�)��QՓ(�fk�9���O�0AŘM�~#����W�?Α&� ���Lw1�Q�M���9q��_ޱL��"� ��4�x�"�ק_d`P�����?����ȑi�o�#5�X;K{U�뾺D�a֡@���qg�������J3���H崑�kt���?r_v�I�+��bdzc<�K��.di��e��arKjިaf����ӷ3�b:�!�6�>Ww����{�H1��Z[!�0�0~�[�}lvh�u&�����b  ���~����#�$͹t����e�
�t�uRR���K/�9|Ǎ������)�����|y<O�c5�tx��s KL��-�uW�u��J�a�W.��d���*�����tɝ~�����s��ˎ�~?��q#;�cP��
�Z�|�ژ
n{�Y�%�R�%�x|�2������\���kMp)��7�����d�i�P_��W���K�6�8�d7�=�A�d��Pg�[���)�H�}C�1Y�W0��/�,���������H8E9�0�vK�L�2��!�5��sG�0⧪^�t���QvZ�� �*�b˅��@jD��0��+������R<�F�k�W�^]��gmȶ4���.�R�T}0�΃7'��2I�/�r����UwL$3WhseP#���'��7aχ5[��U �r��1��9	κ�f��n$"�׹�h��br]Q.���,���#����#!���M���G����"p2Y���ж$w�`Y��D6��u�p�~���lo��S�R*��:E.*d��� �"Uܽ%*S�ۀ �~P~�P9����z�a����K�Q��Ψ����$M���?����sZ���z�Kރ��X8	=%
��;�j)t![���ߊ�Q��D����@ٌv2QV${��*��S�RI�t�v�q��'��Md�B�"�'?�b��<���&W�r3D�'.8+�m�|9�>��ZrF�O�K�0�ӓ<]�A��aa�`�)��h6�<���	�@p�~2v���|> ��v�+8я}52�N�'ڝ��<Q�n�-}ݜ0JA!Mۦs����x�b5ׁ������ڞ�,�y��X�!�s)�Cg6���5'|�H�#ʓM:���TgP��e��p��x@U}���o�g �=�aMo�P��A��x�o�R��S�GL�]�H����C����L���_l��z���,�9<��Y�6̹�O{�su9�B��(K(NKmСMw�yX����F=j&X0c�n�d�  3�s�]��/c�+��fp݄8(ۏ:�$7���J�ܘ\|J���WdX�KG��X��C�sCq�?�oF\��/���_����9 ��;P�>�>NI�jU��r��U~��~E��Z�{j�ҒM&�ύ{�1;�'�����E��7���G���>��5��ITi���Y��2� �94�w4����F@��W9�5��X��ȣ/��ڦT��
_�C"$�Y�/�j+b�(�	�G�,E`r���k!���A8E�J��\(|�zWG��1HX[�mI �sZ�1��[x��h�rA>7P�?|���`v�u�!�c��g�!��N࿂=�ҧ��3�-K�E4$��+P]��sj��h�D�l�t�!u$����R��/�L��##����.��lR�7��NJ���I�	pe�;<'YyJ�i���n,�6��҄����L�/n�5�dT��:tD~����|�ւ�}6�����2���YWF �(�}��k�.�P�X^�SkAg�i�Ћ'M���Q�Ì�}�Q�5Q s��b�sb���D��x-et,��*ڑ,cgH�Ё�'��$��H˞s��<�R!u�����D��.����a���L�ו�B����o��ےυ*��a�-�m/��#���@���=���!�5^�Aj	��k��+�/*�. �;��K���� s�:��P�M�T��!�����y���e�9����us_�q��b�\��_	��lq�G&�5�������gmҔr�Z��s�h���l�X�QзEi�74����\���z���ĝ�<r|2L�q�t�fU.Q1Y����V�Ve��}��1(��=|��=�V��]sj����H\ҧ�t�E��z����w�D����)lGܠ�N����Zr[)�ů�����w�
�pW�r�G��.[�q�h�"�j��^=9����o:�;F�-s��[��U��M!�Z��@e:D�m.T~���/v'Y��b}ئl�$X�9���^�^R��� �7JXdzE�M��^�d���?1ω$�� T��� D���N�X�Ssܫ��*�<�É+�.�C�XT��i�8t�8<#� ܾQ@�~B�G� �R�W��5[�d	Ȳ)TjOQ�v;����;�g�����B��N-���|�ptS_��pM���Sۊ�髧	P���2�����s���b����8	�*��AP��v�2��,f��{�_���i�A�B�[�N�
Q�̳R���[�vA?��"ļ�~�"��G��ʮ���u��]��fp��E��J�L���l�)[��,ݏk>s3b���`�<tɱ����!�[���~w��И�����{~�TX���t��yͺ�tj�MB��l$�"ϮpoT��b�N�le�;pY$M��K���~�PH�E�!����,��*�';��d؟��uM�Ӟs��U�O�{��c�a`�b
Gru���@*oЍS�۴����u����dkO�\�w��c�~�k�r�2b��t֕{��|�?�(��5k,h����w	�o?��AV2��yod��Tb�p�|�K��&CIL��(������Q�	E�Y��y���B�|�5����z�ܩ5�<�߳σћ��ȑg�!�\E�.e��U$�P�k���	����U�������'�}�u�r0}�S7��fm�)�w�1��I��ɊP���_�,�ԀA�:5e�&b�T%"��]�̤F.��y�����.��
 D�Y���P�>�F0;臬ם�4_A�P		� ����Z(7cC�Hi(] �8��g�դ�QOIF���rQ3��0i�Q����6EJ�,&4� �,z���Wc�V�8��lr���~����nͣ���i_#��I{v��W����B�جW���{��OE#��M����9Y�TA�9l ��V6(���z���!f��+=����uh�n�S<�O���[��R��0�Q�:���m���;�7�@�*��-"�`��V�,]�������A�З�l��{pF���B]'�"�Y�<Qc��%����:�օ��QpjȭNX���L���<:�-��G�~!�"Hg���\�]!�s��d`�1sJb���u-��C��<�p���� T%	�+�6\}�Jt�+.��>w��-�5-���5��p�W/hJ��C�[��x��{�;z�����N�6E�d,���/w��J�u��-�f��R,(t�bC���(�?��	��c�˅7��B�p܈}�)�_�	ZmQj5k-����4��fc�|�z�gHK�88����`��6IK뛇߃��e��++6⏍L�R)B�Օ�,�WT�v�߳�?�H����)5�fG75��w�;��Y���8�!t�:E0�y.�6˩�x����v_��t�%�W���������ږ��xb>��n�����`�O�<��:�*=�r� $i67mC���01�M�ӷ~��$�|`?˘P����=S��n9��%s"5��}����iaw.���ya�+� MB�5m�h.�� �9�G.��p�b�r���0����g)�۞/AN��օy��\��tg�'Ȅ/��󅝼T�y�Y�5R�҈��h�\�PW��x�N�v>�]Շ�;	��>�WAwZi����~�\�n�����v�l�����1���_�����!@>����j�Iw�2�h�DXZas�,a�����%���D�~��wt�ed�6��1\�p�����mt��SZ7��'	�34�#a�qIZ/Cm7>��s��I;���+vI����T�	�V�J�:��nc�s���v����;wTǱ��'$k&"�h��ۮS��[�E�[N�k�$VF�G4�n����Q�$�"�ӫ~RF�1Y{I/������ö�"�3R��0?d���.>אP=|�
J�m�K���B��N7�lD�sp�Ơ"S��u�r�K����r>�a�W:��y�
����?���l17����S���U���O|��[>+=�1A'wx�HR�^E3��It�&�R�uQ�NF��0Õ�pu�Q�u��W��H$j��m�Ƌ��Y�c��@� �ń�\
!���_��6����u>"W�puJQ�3����Vr}�3ŀ�0�����q�@=)r'r�Zy�]r
�ۉ�0��g�z��@S��TQ�Y�AP�cR1QLCL�T%�ym��xЗ'�Еb�ځ1�$j�\g5���QY�u-���`4`è�0�][Uy!V����Ϲ���ז*(�Y�6��d��c�R�?��S��n	����L�QC����c��B�_"���5��ef�H�t�U�{)�~��k�yn��L�b�!����R�.G�1��}�PM�H"��Z�&^��?3z�����霈� +�g�ͩ�;�d!�ɟa<��w�veڭ����k��g��`�R;�5�^�-6�O��F��~����wf@	38��s��b3�%�b{�)e2Xۜ�K�nG��@-��d���WG�T�A)/yl�%��c?i����I�}����٣[�;�X�oYcDj��7 ]��%N3�>x�oT�AZ��E�O�CkO�4���Uw!����3 ,vI���nMn"��h�@?:�� eU��x�цّiF�-<׾�EE�l\*��A;��$��r���-��j3�M]�;z����<�UDӑ������_
��>�ݢ,�:�\����MO1���:Lz�KZ-ip�C�(�3Uoh9�m@Ulx׆)�z�z� �>�,6�c��g�ݍ�g���b��$zr�6P��&��P����'�Y	�N��=Sa��)�0� {6���:#U��$�:�Ǎ��`,�?h��(v�р
)�Dݴ�aX��H����X�����r_5�w*RP;c 1��m�M���qR��L���E �WǴo_b�3���A̐�Aۧ	|��DLD48����*�@���7cY�!]%�n7 @��C�X��{=v�(^�HE7���>��w���ң�Wp�3.��=���p�Uט�*��T����`��~ޟ�e6�kϨ	g�����K]��n�5�t!Wb�>�����<�
쾳Z�QJ��f�}"
��K:n���-�7a���{IQ�����G�6���G�N�Ռ��-�{�1

��a���m�t�>�0��%�a����#�&��s*b��Z"?�iB��fL	��kܫ�}� T�f�a0I�(�0�x��.�h^���J����;j�"�W����W*����D��8��{+���^�`�L]���f�P��$������V��K4u���%:U:��)�Δ��C��L]t&:�h�k!�|�3E�z/|1�m�k�D�G��h���)i-��;-�27�uz;¶�L���QR;��hH'�<���r}���8
�o�7W��qr{#L�V�|a8�<>��N�����g�/���,s
�Y�W7)m^�����'jۮ�y���u^u=����m^H�I���?��?�E���:���i_��"5}��!�M�����WBڊ���4mѲ�����*f�Ɯ
)��Cd ��k��u�A{����_rTa����I~�dH��.�n��#�+� 6*iD4U�|��p�F����L�%��Mئ���/��I~@�/�����=�;,�(���Qy�z���K�m��T�c[7FN���wH�������Ӓ6���8���/b�ڊ�QM^�b��AQ���Y�&�*�N���FI��"�rS�Je�f'�sd<�PJ}햅K�x5�kd%B�EJ�6�=v)�Uh!�V3�� �X23�2v������;��}>ߪ}27���i��� 'WD���~���z-:�a'�~@� |�U[0��mo��)'݀�9.r�'��Թ��'��dъ�W�ed����z^�طM��?�u1�c�W���'gɺ�v�n�r�ׄ��g@\�/?�ݏc�8��E���k�����^#vV)[ʑ>�`8� <��y1�P�i�m��]���/B�4q:ZY#�$����.��	���]E�-�cIU�������)w��R��#:��Xl��w
�?�/Vo� ��:�[�'�ϙ��@�Tz����b��i���[vr����e:�~b@��:���DP:&��g� �[���ߌ�K�Sl�$�T���ŝ��(c��=�|Z�̏F-)E�JJ�6>G+�-{�4�n�����j?Rj���R�I:�� �o6?��Z���[_\�Ws�y�vOX@a��;�%����z�����R<4z�ŝ?E�"���Vϸ;T��=����J.Yɾ�[������ۺ�"R,���1ӬCN�}�½�����tI�
E�F��֭�6�[R� υ~����vS���Q?�XD)����`<Xǈ�;����B7H���[�n�{�0���\lh����ð���t@(�
�=�l�H��/U���y9�@�
ڀ�`��f�B�Z �=�mT-��0N���8���ۡ�D+�4@���t�w�w<�ßj68�?��f{Y�6礐tiA�dE��uN����XtBQ��x �G��1I��TN�閴��#���l�K���P��ahz>�Y\�z�˧L�9���A�����QE���p�y��<[�Z��Ze&�\�'n�ue��;����A���o��mrq|���r��"F������������z���K��D�w��X�9���W,7�\�+�$�)�6��ƣ���%��`�ls�s9Kq�����%�d �
�%�F
�Bl?l3T�Z"V�bڢ�|r��9�9%ouu�gVoQ�뜒��������5�5�سa�e�0G�ߺ[� ��%�9�h��G����`������خ�Dz\���L���T�]ՔS�dx�d���
�!✿ۧ&.��������R=~{�a%��fJ��6e���T��ǉK�`�T��x�/����0��s)�i�+l���.�5�c�[J�}���L/<�E�v>��?�l�JD0w�*�1�f��F��!o{���v��qCf}l��Omz_j~��h:(�֩�����"��궬74�lЃ��ڞ�wy�k� ���rc!c͢Ih~9^��	Rt�Rr�x��>������� U���;t��6L�� ��K~SeP
����ia(���^u����}���k3:hq���>�0L��
ogO�5��[R��X�Z�d1�������}c�N�KH����N-B��ط� �<�̣T�������d�h��+{��+��6�+@���	��e��!Sq-��Ʋ��%��mi��q@���V� ��d�>֪�tEx�{��L�v����AM�8Z��׾��r���cݪB���FD��c���Q?�!ȸz �/��m`�!MG��e;`4)��CZ�u^�?�\��b?n��-
��l��_ ��yS��H����9C(UD�ؚp#�%�]][D!�d#����r�??��%hUJ�%	����f���=>�_CHF��b�Ğp�x�-.V�� \;x�j ��"����ɂ]�3=&�Zy��'L5���Qh`�T�A@����G�(?j�0�Bf��d`t��":�h��R��w��ѻ�6.Qr�N�W�\[���P��s�h�����1�dmr�IΖ�J�|�ҏ��!c��f�A�<�����v�M!���:��E������hﭭ��O��kJ�n�է[���
�ʳǵ�ݵ𡈵R/����x��S o�n��l����%�8��g�M):�{��N�s��Ӭ=u~'�Q�Q��"S��˿+F����[Rmr%T�.5O_v.\&��J\�����c �H�
�X���d��:�͚�ݙpn�"�X�����1^�N���z��	2�2H�ӄ���+z�P�2]��KMu ��sf(��kj=���h� �ɋ�[o]`�Z��+"�vFP��
B���Co��dc�d�dj���Mc��W�1
Q�m�@[+8�� dā5T���f�}srh��)����WO︵����?	�8`z(Y��I�//'�����`V
���o��.����	ˑ��A��E�F��BKo&������\���&1�i�X5Xf%{މ `�S�WG76d�Q�݀�m��D�'fD\5	����Aڐ�Iӭ���rnCg�{�������4S��fm|)�r;�~�!�ڊah�d9����ȸ5=
�b{�K���G���[r9�3c&_A���4��J@�u��XZC��?l�;��hx�'�5�U"eCy��hc�+��f��;��Ʀ@��׫)A� ɉ�=~Q3���`l��N���q�6������Ps_�/�2��;�h,�)�w�;� ����˦��~������z��2a�)�7��t����>E�P>.]@N�I8M0��xf]���t<��`G{G��XlxV64EB    2c82     9d0ЭQ���B�1|��IQ��K�n/g&�1�;C�!TD�᲋o�x�L(ނ��GA�%�|�?�g�,�$0t�fS��{c;׶�?&I#>�7��_y�?�L�7�� �?A�<�B6 ��j++Mу�6w���v���
,�ט9#i!!� �F�x��Ѡ�����ri��F�������}��0�2�u�~܊��s�N�?��)�P��F�	t/q�Ʉ��yf���bb�=+�R�nn�+��0��V�@���,�ö���zi�$|�ڗ�Nok̂�&u�(Y~��Y)��Km-)��h�����P���^�6cH��ß�ҵ��p$���K�����܉_��Q�Ьb�ixU�@Hd
�蝏H=�捻���.M>��ߩ������֟z����ɽ��Ѽ�\&t8��0j/����C;J?I]��3���S��oJܕ���_�{�$�҅$����.#{(�� f�������������q�2�I�<f�X�AQ+�zYYtޜ�{�b�lW7����Բ�i�Ch�4��=�	Q���2DX�JLQ"��y-����>�p�n��Ƶ#��(�	��ɈbH��~�wcp�hH��&�n�Ayݑ��4�
�V���B�uM�iPĞ�k�e���z�E��o����A� �O�ì�w���������c�/݇ν�Q3N�W��9nD��x3ù[S)?�#�u�n��9"�#����9�
oK~�J����#�����Rt���^7-z��4�u��f����qvf�s�+�=�}y7;I��2l����LdYg�8�
���̶�H�%|:U�
Ҥ �rU�]��p��<��i�p�۩H#q�zR��:��L�uϋ�~/���5 �Z~O;�Z7c�V�_Y��Bb*�|;��(�V*h��Ar(��Z<���*~���	�07��ߵ���kX3=y�{;�.~#����օ�6���)�U�դ1ҏ@���n_����	 ��I�d~rxI������$��K��x��&�}P[�oL&*i����<K�S���[Y߽TE�1���� Pߧ��hn��ߦ�*܉��P�ZÑ��9�[��s>��r��)�j��p���(�+��R'�K�����AL߶w�g�**C�V��Ɍ�Ȥ�x�8$)�r_�\$�t�"j���9��AY۫,>f�l4G��+I}�	�#�>2����I-�Bѯ�n�V���t�Y@R�(����喫h/d+�},f!9�6/=��a���=<F����j($緳v�W�~- �YD�Ή���߾n�qU:����d��O� C/>aK_	rqf$SJ�K�m���ӵ�a���0	!3�t�#�$�)ї�%P����w��9��.�Jo=Z�����~� �&�B��d��&��>t�C�w#�h�Bm�*�,u����=M.�A��-$6�׭Ϧ�p�D��8
�T���]Z8��S��DI�`Z���m�ie��s��{�y'�3`,=L���8G(�	��)�:�����ʎ�};|cl�,)����b4����8ǻL�5I��R�D��1h�N1�~`��x�(W��o�{���ӕ�H�
 ���KK��B�����:�>�"�]P.d������g�ܙ���Q�Y�@Nf�fa^����T�%��������9��e�Fn)��
ir�纄�0,�'1zڤ���wlKn�u��#+������P�4����!��� �z�Ȧ(���h`�Su~����y��k�l�@!u�3'{����L�d��B���#l�BI�t��h>�\l�1�4HhF�^ {�X�g��J�!��d�'�U	�S���B3V�-�Y&_='^���+��3p@�.���G|P�"�>�Q1�f�Z�GT@T�p���g���9���-<�P���� N�5Q�c�J7�1�e�ӓ�w��Ksr�	X� fu:g��A��m�IN�����uGT3(A��mj��pS��Y��!��.{ЌR�Ґ./p^Wt�fD�Wf��joUYˬ=�6�}���P��Y*��%���?�'൫w�=�2����kV;�׻߱`�B��8�C��d��J�$~�\���Ӵ�߲�V��&!y��@%%�B�[���1Š�n�������������Bɦ�:Q�e�����8�65ʞ!k�Q �et�*�V�EO�]7�"O�L#ϧ����dȵf��ˠ���4�m�mÃ鑩����6|,�#�����h�œ�$Y��ˍ�pi+��F]��6y���1�c&J<�f���Ț7|�Y~l�#7\��I��$�0��$�ٝX�%^��M�v�=�Ia��-F�	�+�M�3_��5���;���\y=���rx�W��M�~��D�a��r�buQA*RP>�b���)�TN1�]��#x�B�i�,���#@2
>����V��.�[է}�6tA�� ��qm ��\2�#��|�