XlxV64EB    1573     870C?�3��D�)Em,����%�釣�-n�CR��q�4��1S���()' Ϯ�fU�O#�m}�����.�[����o������|j�<l>>�L6��xpo�!�DН�Ou�6t��ލ,n��������qlDdR#����7�T���7�����:0ݼT�E�]�s�%\L��@U���g,�j����Y*X��P��ϴ�&����O�>��+���;S�§�����a9&���]O�\x
	�5ۘ��ef<Y-�y'R�J��^���^�$�~���R�ah�ރ�~�,�eF{���B��y�j��X��Lk!�
S�/�����9u���q¥a8l\���!9��<6�}[�CY!I�U��$�p~�vC�s����2�Պp���vBTdxKBr˵a�t�3���T�`[��,��%�5Tu�u�҄[�
O��i��1��k #]�\yݎ�L5MQ+n[�ԭ(���7rn��Yh \���-�*t�Պ��+�')�$�!d�"������Dag���9�BJ�0	�үbt<R�_�9P�CBou��"O㌌�^[^H��Y�j	1;쪘�6>��Aj� @��� y]g���Hъ�������O�cLo�8�����>�2n_�wOL3^����f ��A�z>)0�]B[��tr�|�M��Tz`=�t�]A��
�����U�o����D�vv�:ک��]�^X37KV�ή6�D�=+r-񮜇'��f��`�����*���yNMh� _�2��(�1�X� R&bS�f|	���@2�e邷�7�]�f�C4? �7P�s	:P�茊�r�Uj�lqbk�i"��+ڳ1ʳrV�������%��c[溞���� ��IH�7�Ȉ7���o�I('S�gs�.�%�B$ ��1E�0R���U��w.�C1�#ʅ����։/��ߐ@Yt�ɬ--��ҍI�|�C��q������w�5�\G���U��?�h�*[N
�/��4�*���R_qSWDM�ƹ8�L&|W^�1>;b���2�P^����yr���&����Ջ���)#�Y#& ��˧>�/z�+G��Q��b(�ҷ�#V�_/54'|�ضv�&��{����vt�N��t�ޖ��2%�d���Ω6�f�L�դK�g���u�{}xb-ɼ�x��t�~��c���cf��jݕ��(�lG�<�X��Z>b���[ �Ew�6��:B/�0V�!�d���V�\;����X�W}�G���82zɡ݄{О�~6�Dt�1$8b,Ss>�12�ЇϬP��8��m`ӻ���N���̷��[�Ix2�*�/&�E�y� �k��M����_����
��r�ZF�Dm���Y7Zd~��˸��u7Y�o+���AN�6��Y�Rvё.6���9��`��E9SJr��
���W)���3��5�v�	{��XY"�Hk��{ϗD
b\{Sr�������g�d���ˌ�+V�d��$7&'ʸ#]lz\4�/��nmv}�b�~�<�Z�C��5��A,+sMY�I�~r	\����vJ�+vE���s��!.f��6��b�y���g�=��3�A��L��*���{�qg�y�j~����?���/#�1�8fXЦ��d�I�j�8�2��(}��O\�U������0�� 	h��@-�A��3q|��%يEi
�yH̡�~h���r�{���(t�l�cl3�w�����=Cº&�TI�a�R���R�U9���Ҷ�1��FF��uuzF�\�nc�P-x� W��oe�&2zE�v���͸cߢp��l�P���@�U�	:��8����7(�M;JW%d�h梽RoR؝�G� �bw��O]P�#��5��ŵ��� Z�z�k�E�f��A/h��Nv<�ީqf�t	��F��7���;VTB�����ne��җ�nDA��q�A]��׿�����{g/o�ߖ��lN��� ���'�Gblj�l�/�������}��|�J�Q)�;� �g�Ȭ�D�����g�-�!�m�#8������m��{���7aBT���xlG�Au\���f�V=���8h���lH.��ܛ�l^x��r!��G�@y`��� M��'�����