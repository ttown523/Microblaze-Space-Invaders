XlxV64EB    fa00    1ec0�:���@a�0����b�x�h�>}y�|�M�4����|�A�i�2� �����,���CfA�&ÅS�+�|����6���vU�q�a\EM�3�`�DtP�O����n�hB!���\���p�"J�v8R��;^��  v;-�ƚvĲ��=MJ2(}�.v�B7�C
~a(��mK
;.�O�k[��m�?���P5�Ů�u��'Y�m�����p���.)),/�&ި�1�
m�z�S�3��jPC�\%M�/���(o�4�~T�Qe$v�۱��B����>ڑ�G�lc�X�nS
ǰ�C}�S#̛���{��ޤm=\�&[��Z3��ԹT��'�. ǃn�Tg/c"�t�ζ�k��H���x6�Z�ѱ�����K�D�N�K�D?+H4˅L3
�4���5q'`%���1[�n+�t��Z������Du6��5��'[5�e�:��,��"�V=����h+�d����Dc��iш)Ep�r1����Z���-Gw���y�twjc��[�R���Pap.�˘����\�1�%䆨k��q� Qҧ)���3f$$��.��עgJ0X�h����Hc�ݳQ�`e�{(BOAY��尯�K�̧ߠ��$q����gc+ZgI�<����Fv����]y��zT#��k�ҔLd��ý���7�q�/x�:uN�u��n0l[���n)���8���;:f�x����j�4B|��"8�%&�<إ�G��o����X�E{��v���O$x��d����/_J���R�m؇���X���0����So��p����j������#C}K�-�x�݀���0豨D�E�Rt�w~�W����c8JRi�h�r/���Q�ތu�����Z���Z|���ܵ�*/��F�U	�l)p�߃���3)s�����F��B�84�~�cJHN�v}y�L���	}�l�"�(m�}c7�d�>��A#��7_���Z�|��m�2�&�d �|��+����ؕ���yU6!���)5\���cn'���f���q�j���� `=70B�j�.�:Wb>¦��!"�NPs�\�����������m���`,������dͼ�(��Ʊ7Rv�\>b����Q<O��v��u���q]u��F�#Vs%�L<�G_}��:�R�S�5�R{�N��f%�����V��rkc�L���p�b�uA1C���$*�gp��Ht��h.��/(�Ǥ�g��q��� z2n����O+�Q���5+���Y %*E�(�� {�$�LGt0Ӣ�Qt#���M)�=|���t�T�K�� �엶P.�@F.�ݱ��$��l���獕~��h�Ѧd��z���Ԏ�t�C�`|�N"�p�E�G1Ƃ��l� �
�x�,��ĩ�[(q��V���ad����X�
�TȎQ&&������@������-���gx	ـ�W�?�4���� �Vc��"�9Hl��4ϟL�Z�Q-����,��Bknf�Q�m��ʾnzo5ι���,Ny�?'*Z{��ʓ�H���|�4��i|^6DG�Y[�a�����M� ��F�8}E��9�Apfە%N8�?u�mqT��c�?u2�z���5� c\��Y�J�9�؂,s�6]8j��^�#�z�����-we���|�;�/��h֫h'�ΐ���z��u���ra�?�-w�����	\�_�����ˁD��,�h;��++�����,�/5�X��ά�J��$D��6H"ΕRi��Ӯ�9��������lV���F_@�����Qc��a �o�՜��Wg�n_��;� ���SE�D�Fͮ	bԺ���^靧r��� � ����%q�'�S�qƨ��ժ5%êk1����x��=G�O���YR�=1�bm�U��BO7}
�Ψ}�UÐ�+�G�0Z�H��`}V0�@&�����Q�$��4t�]��M�aw<��3��NC�ѹ�зZ���DA{dJ_�m�%_U[nD���n|:/������t�Fbk%��;�HŔzD����ZcI�hA��� �ɫX��~z��𷈒h�)�J�gD�t�@�id��'ӟ�ds���i�6�9��%@cP8V)���V�*�}m 8(PO[��#jCY�*3jO<<f
ygH�J���\&�*N.z_'p�
վF-Wt���?Q��r!��E���*ϰ�'��ہ�ob�r���2�T�T��	 ��օ�O��f�4���=��;��p��6�Y0�"�o��oR^ ~��AIh��;Ȕ,����A0��9�������q���ZS��� A!��. xv����cU��|ְmo��,�RL *���d����9&�[��%�BH��υ�[n�j��~��*4b��!qA2���(I�l�Z��P���΄��tp�>�賱5��Ǡ1�3�3f�L���O��R��˨�L�;pE� >Y�F�_��I�w��1rU+�zn�F��b�;7lp�63v���ވ}ѪU@�C�@�L���Zęgq	n)���=��Ry�/Zd�i�|������..K�yv>r~dͬ�w��4�ԷكG�	�v��^`c{X!�!�L� w�٥hr���+T�o�9�W৩�"�S=����[cs��c졎�M���XQ��F� #K�wN+Ec�I�RP��KG�qִ�^�Dm�A���۸�VgG#�S�Ք5a1�y�=����ive�.?3x�^���3L�¹y&�j$0�X$�e��C"�o��<�l.�����E |a����.��r����R~�	���F��ml�0&���p�K4����������dhQ�#�������{,�Ƒ�ލ���Z����(uWW�ּ",ϲ��꯶�� �a_�*u7>�C6d]l�� ���C��j�Ob\�:
|��C�^�We���D \aj�шV��ꖌ�K㥛�����j�4i޾���N�����"�p#��Z
x$i��u�����A;�'g��쵩�rUi��E���Y���m���#�ea��I� m���]��{V�~��	@(Y�g��H�ӌ����m�޽DU����)�L�J%W=�C�6���H�H#h&\�b�ȑF���,�;8H�hS<����{٬5���K]���qh2~g�0����>2��{�+���@V��<		L_�R;Mҫ-���Δ��7���N�u<��,NA* �ɚ�}2�J0�n�:��;<�g�kj1�Q����ا�>k�xHȅ���bʮ�_ZS}��B.&��>�f�0�
rZ�=���+�#�W�����D�VzyD� �����z�(�����f�ḍ5c� ��B_J>��.�N*f'��fE��
� \�2�j�8���]�g��/�������'	h0|��B�|�b�S�i8�	��e:z$֞l(���nگ�W*�W�D�έ+�Ԓpf���󏕚1|XoC���9�e�&��a2��2�x�D��"5"���7��ۀ� 90�=�f�Y�i l��TԈ�d?D���Tv�J�"���:c4m"�$�]O��-���EŊ2��ʎU��MS-�Gp9�(J�����38lQ�!�,�O
�=t^u'E�'����9�IO��M�Ҕn1���,�^$�պ��ΐA���僜8N�Qi;�;���35!��tǡ�X�Ɩ�z�2���@E��d���Uq^r<�!�N�Ue�����z ���4��F۬'1ɤ�\� ��^&�KA(�q�q���
�]�d3�`fPI�0x��r�-)�rfك���4�ttٓ(�u1�h��f��^C����9�<w�w�N���~��=v[��\�M�a�~�ڑ���#�@ygi�iᴔ
�0q�fU�[ڪ������H<�&�n�����/S)�^$�u�Ր�;�T�K����.PM���|I1e����.�ޒ��"���)�����nş�r3Q}��u`�^j,K{�}RCd��lh��`5����Q�@LRd1
Ο3���+�_��xHl-��^.l�O�T2��m{֒U������]h"��K��֋��7�������kkxA��z�:���|m?��/�w��3;ʹ�&@�Ge]��/� �6���I ��-[��+�d4�O{𭑁MI��C�`��fy%�tmc3g+_�ʃ�S�-._��ǜ8���3��%Eu��"���X�3�'��Q*V?��� �ٽ-�]���a��{k�%-b�l*mI���qf"��k�=$Q��hU$����So���m�GP�&qϝ^x;��O��Y�3�a(�B�ס�d�(}o��}.Ld5�i���Q���e�O�b���6�$C��U����+) ��-܌����<C��П�o<�ƅ�s�6rۀ�L��X�8�'F�$��K�k�t��	��փ�G*�2�4�b�����P'm�L##"zW9�=�Գ����K�M&
�N�C�w����ɇӱ��؛gf��q��t���,�U���>��$��n������+�%<��Y<�@�]Ǣ`�eu��^�������~���𮒟���Q�&:��1�2� ��6^
��3�oMc�7����@��/��1T���Y%����@س�ט�~�����ɹ�)���c �n��f���8�r ��:�5ؤoJ&18��]��4��V�����r�x�kT [86�i���:�w�W�w��
ٍnW�x#KB�HO� �_wl`�*L!�� �S�J|�W�A���x�����,���Y3#eϝ���h!�:�}U	=���1���n{F�V��CX8͐/v��L��;�%}��Z��&�v�,��bD~��#��RRe�^<���cx�=n�>�z���Ґ���Q�2��(k�d��eNCy���P�b��9��_h�t�!�Fs�?��$	ڟ��!�n
aTv������9�UܼKJ�v��p�;��a{����3F� �EL���dµևs��PNy]q�pAM(�¸�4�wV�Ab�m��載��<���?6R�r�`�z��1�?���F�U����'��	��x�vy?�l�O[�
�!x���Mm�������b�vcݾ�kK
�d5�u���屶ͨ�fq۱wj�s� "	:]H�meP���R��2)u�7�v��/#7�TA�Rds��iV	����|c!�S&�X"y}i	��K�	KK4['d`LT��[UQhL� �WA*#\T�2i����)�x ʘ|v�\Qe�m7�K�ZX�"�P��I�|�t�f�7�����.A�Td���T���7^���,���K����	�������z�5ms����5�Y�Au=�46g�W�,�O����7?�4�
���j�j�O�Њ(��K�����=!��e�a�X���5V	�x+���ݽ@���]3�� �@P���!���,�"A�|e�G������#�'t�[.�x"���5Ej� l!L��͜R^'�Hh��b0�a�B��}��r^��<�TO=n�V�j�e|^����'h�YMzs�4��[#ʑ�x�-x�g�|��+_I��3��˼)^����\P��]0�Q�h�9��ө\���o3[����hFn�Rɵ2	��@a��
�",�ߍ�C�՝���F�o��Mk��t2��|��CZ�4Z���v�劵��,no�1!��6�Q�v�rZƳӅQ{H��O�&�'	� qŵ隽D0����	�"��MQZ�ZnRMJNQ�8�����Ģ�BZ�A�����(36�XO��C;����|q'?7Hʶ��q�@�bxg:]��q<��<x���������� �~��}+rN��I���w��#P ������qy%��#�)�u�.ɓQ�����"���E8j����8l���hqU������߯}�;�fy1�z���*O�OW/%P������ �/3��~����S7��gX5�YS��lU� �XLY�m=[=����V�ɛzAjS��	1T?$~����	�h<�d������s��YB�A�,݃��s��N�hZ@��[�E z���
B�Ѽ�#BY�$��^[�Lŷwt��$�ٙ���Ft� �*F��v�tLw�� -k\� ��$�~d�L������v���#29ϐ�"?L�y���9�������v��3��!�p�V��	eۧ�����Ts���́��E�O*q]�_�K8��n���V���Q��n����GN"ףm��~���]�Z��*��b �^xA���D���I+�Z�Xe�d���3�kHg-�u��/�o �� �}[�9���p.��,P�e�#�v�;|���A]!��-��4�٬�]��ž�0���~���Z�+ֿˊ�m�-�W�0j��U�����D���PZb�'96p��g���
���JVc�)5�m�����Û���R�c�#���� ��ٹm����<���s��>�R &�`�B����"�\GXs�}a+w�H�e[�VY2�a*ۚ�W�� ��D��(���A�s��5kj5|hh��4��U�&��?�w�+7�p�y�vj��y!� =XR2��bÃ'�����L[�zLR: ��V'6�["���K|ت<[?{�_`V����q�� L
-���7���o��͐
Ĳ�D���0k�A�n7l�cT��
aæ�f/����m��r�wO��|��t��n#e�9:[���������t�AZޠ.����޺E�y�4�_�*|ōm�=���B�孱.���t�u��V����U�֍��Hw�ZǓ���	���%T`����{j�6)�m5.��S�x�=���i���Ti���Z�x�%(�װ7�,�gp�;�������.��;�[Jl,P�1l7X �B^����똊֟���1թT�Ը��>3�DK������t.v5E;�=c�q��[�����TOj�ɥ�4?QCt����7TI�S5x�Sa�6k��s��A�$�VD���D��F���O���%)=4�+��F�H�hG(��)+�Q�%.����Q�l�S#|>
i<�᧜���\������'��G1W|Hܰ��{��pNi�(����&�G3i���H#q�W�%�Bo���E����z*.���gU��o�����ǝ�����S�@F%c��l�k��D���[9�k�#�ͺo糟�F{�Xj���|��ڹ�߭�)�v�Hj��q���Ǟ�%��t��"�	ݢ*eT/M��M���)����4�W���0�L⧱�*�9��q-y����es��V�S��	���Cʙ�*y#��)Z&�����h^�i/�2�i��8w����rd	וq"���vO�)��ӵp�`�3�E�`_�V� �|;�#��+���/c��l��	c�K��M�x��S��I�gJ�+���\�������Tn:@G�b<[�J/`-|!����u2Ɩ �����W��	hcoC�G (;�z� �(F�2ט��-,�cTv��qmyL	��y�]��Ꚉqt��tc�2cb��t���`ݑ'��_p̠�ѕ/����v�	�mn�יX�]��c� �
vE�6��!'mW��F��X�F�Ѩ(���7�">�7�j�e"H���'�[���:��0>�-/΢e�n$�T9�L瞁�U����|$��A�[G�X����\"E�XlxV64EB    7be7     cf0�:��VT�+星���"�K�P�������4a�������W��Hj���_TPt�>!]�B�z��n�w�22 �@�{1s�1<�#�����l,�p��&Y9�_�f�2K<�J̄�H�M�3D�+�ӭ)�댋��,i�8yo(v.�_[���+eg��B���a�"��r-g^HK�?�e��%4q
}���}d�|�)����8؟C1V�ː{^&�hD�v�-�?��Z�>FA�2bO�'6< �У�^R�����o+؁Krw��	�Q�Ƙ��	�1'Xάe[�2�K<� %�!�p�p5]m��܃�4�7��ؼ�+��:��Cj!^r�����	X�ɂ�O��ZK�nǠ�p�&ۏx�pK��OJ����O��B ���?=8.���4gL�k�Q��0
3�i$�3����j�C�6C�^fK�CM���Z-"fqC�1Bt�q*�J���zb��m;��l�,۹�M�����R�c�~��)pj Z�&�&?֟�/�T�ߤ=3y��-m߯?�be3�ε�\P�h�
�_Q���p b�~XGI#��]���ʝ�h�<j-&�K��̍Ĵ�L#�WJi�@e�@bLmY���I㲤�6л)(V���r��;aC�]n������97(M�ó�}|��W~�����^u�E��G���Z���+��q��	����0��5�K�,V7#�+H�$ts[�}y�B���Q'r)�H�ҵ�>`�����O��f���d����ܗfp�L��qx�7X����]r//�j����~^7�O�D���Q0�S�UV�k���3�z�=MJ��W���s��UfP�N)^q�߄d)�v�|͞ڙ��L�(/�d�-#xQw��q����3(w����,23z,�kFF��t��k�_\�7�0�[�5s�./��ݳ-ǻ�.<��C���Ka��v�9o���7���#̶���/)zz<n�%#$�LS�j5��p�TP��&L5�^�'�0;1�,޴?�dU.�c�V�P�A5�Z�k��/����>aE��������'�ƝMA[Z@W�-�^���rH	p��?�}��V��L`�ܤ�����y��K!�F��ku�t��d���t�'R�7���K��V��ל��t�J��J�'8E��Rk�ΝS�uTZ2����_fD �N�S��nnϵ��͘������Ȉb�ZڅK�$��_3�;���f2�$����+B+m����4���s���+2{G&���a�x���Jt��E�q��An�jc�-[�#��~�*j���	�|kP�N�Ah��͘j5���(NZe�aR�vQªr����w�/z�S3sv΂�-�Z�cR��q�MV\��;R����,�˭��vM���wǘ�Vyg��	��f����?_Y���`,QW}T'�л�>��(�3�sC�����3�����m�up�x��4��w�{!uS��>��o�t.
!�D*����9Z�2ʿ��}3p�����F�2�L�@yq�̹'iim��9�����q�qt����}�REd��f��E��m����~�?�����k�	E�ϩ�P�2��l[�:�Q띥T�1�����VU�e�67`q̝ �`������/�x1�N����+���R�	��AEPgW'?�#�wvX3*���bQ�Kd�уi����>̈́
��C�������� bN'} �8N밞	��2ƣ�E��G]ŵ!,�!�A�6Eb7�}���0�_<��%ٲ\1��R1����{oE'޺��tԱ��
L�i�W�����U"M��5�s#���ÿ���
R|���Y����?���[����Y���qo�j�}�z�>�V�f���U�p��S�n���J,��=V@⨁5�A!���5�Щ����R��,J����#P���]�{�׻"ZB�z��x_����ކ�4�Z�d���*�f�9I�.C������x�'ƳF�G8We-r
�����IwL���9�8�<I�_YY�=��j���2�'w���m�G�fBAq����7����#��>�}�k?'��l��`R
��D6#Jm͐�!Zd����`^+1��#4�I�ī� K�)�<�q B|,�=!�+�U׫�j���	�U����M��k��{Ec�����������i7o����Ң�GO bG�Xi�0��нX�!.޸3����֪��U�E��E�����;x�e�������Z�9�&�,�j�3�Թ������mU_B���'�s�O/"1���aD��mCm`ZZQL�'"TaD�����oJl�C=�� J�y~t���P��43�_L�r�.(T��f	����b��8v�/�5����5]Pλ��*��R]��?�]���&��VE�|!'�u��#�#�����7΢�+����O۴/:��,'�X��f�ܩ�h6��qL�����Sy���?���2nxS�lSRֻ*�cp@��T��ùKl��m�T�m#����#��-&Cgo�����_�2�F�e!�Ǹ�[b�o/ b	�*���&�O)�"F+���x" "x�>e�z-��y�j�&A}�;�4��a�g<�6���K0�b����n�6C�LVp_8�
A�nA��Z����N��o���IDx�suϴe�Cc�܊��T2�����^���:���_����ǎ���V����*I����X��*R�=��es�}|D�r��
�UJ�wm�OQ�����S�蘨w��>/�Ńt�H�ZY��kҖ�f0�=���|'q���i�?i��p^t�/�D��~ 
z�W��g05ѽ|�_��T��xo�;*���S�~��K�����G7���-D]Hw���u�Q`�{��}-�R� Lǧ&)m����,iU�?�t�$� �Ôۓ��i<c�x�&+�a���$�'����m�7�5���G������Y�ύ!,���Np��*ཌ�!�z����#��(�@6�U�n�:�.+�� w��$p�2�-�>̆\�Y�K&��n@r����*mHc��	9	�wK�d
�ӂ����ݤ �܅\��B�:���<���7ovƒx K���Ǹ?�~�g]�g�P�[G��58���G�)�a���D�%�<߅�\�r]�s%^�ց?Y��%��,��,�c��Y�{|�ŭW�q;��RSd�vd�#e�h�lp�'(i9ʮ�׏;
w#�i)��K����*� yh��Q>|�;d�V�b�ёPp��r�_�9��(��E�\����h�E���Cją`����KN:���|��LZو"�ؼ��W\���