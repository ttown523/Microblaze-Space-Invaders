XlxV64EB    55ce    13c0T�47��ڿ�����[��/�� ���λ`�X=i�3�5�����=�Pm��gh�i<W ��rC27�Yå��c 8�]�{a6�=������-�L��D���\~.a����,W�%�h�Qb�-��ѱ��g��)�K��a��=ѽ��>.pD��c�Oz���\}��Wd[i/����]f��;�!��걕h���&Z<�nk����t��0x�>�4�s7x�����:�@�����2@��c���&*���ʋ=e�R��o�n;�m.wy�=�e��m~a����Eg��P���UU���i�m����x���,T�_t9�=p�����U�f���D5F��q`���-�Ɉ���ApF9uv�P�^�����g5/JN�r�E~4�!�c����O�?�Q�\:�'�L�~
4�=��D�D�&a��� jkK4�UgR�C�)-��dM�����qI�B��O��S?���86CU��C�w�¸�ثu��R�X���xy�-Eǔ���w"��)a��Z"Z۸�Љ�U�rΊ�{9�a}�O@^N����@�*^�E�~���3��Ԅ"�:wl�FA�O��~����d��՜8_?Y8�\�jC#K(h���6�kn�5��K>JՀՃ��.���0-��
x�� 4.�f/i)�w��hVOW��V����a B���	��׻���w�b T<��4�i�~$�%I��2���H���d?<����;�P�{+�@Fɇ=��� }ŦԤ�'չ��h�EY`j��49w�E�i�z����j�鋹cF��w|�ֈ�l���y�C����)�z��9�j�}�΁ �4�Ķ�{a8F��b���e�u*.���ې�u��-x�ܢ�A1���y�k�GB��B���uEږ������ϊ0��g�oQ6&�o��]���̭/�ϵy���l�����g�$����8sE��D�V����~�����}X:�_�u�Q�S���}�H ��^���H khƸJ�V@r�|>�I���>G�������$g�;��`0��q�c�K)
߹���WG5�Yo�A�_�M��jw�6���me�BY��ʸ�F@�g�&پ���Ǉ�՛�Aă�DXq�H��2���K��Q��<IO�+2}��"\���h(���f����Q):9.m�BH�G���`]}m�荁�Z���������D�#�f�'Ev[_k�벺y9 &�D5� ;Pc �����y6���t8�L�d�S!��u����P�K�O��E+ʙ�u�x����Ny�"���:mX��	~,�~���8!��񕝷�Wߞuzi�)��G<��퐐����J;�8��B�� (c��ST�T��\T| tܙ�B�5i�4�hz#Ҧiln��K߿�.�i*�9��@-U*��T{J�����RY&�<a��1���N�z�R����R�X	�Y�������1�<����1w@#Z�yEnA�PbX�&̴� E��N��	PW[k����Fq��0p�G�Ww\���.�.�ޟ��<�46�����8�v�<�V����g�]Գ&�̎"������I*�Q�Q�+�c���ϕ�1��:w��Bk<r���
��JV%��M'� ��p]6��mm 8G�vDJ���Z-qn,��	`�������yɜ���-TF I'�5�p)0�����Y|��/�A�Cv�ブ0�bU:�I,0mA?��������/�' p���P�Bmd]6�z�2t/0��콙�.X^����9x�
�߸�$�?j�V9>l���o��y�,ld�~>L�wtnڊľ�������qW����h/2�>���M��TH�?����pP�X(!K���{^gHo�+G2)�ix�����'�Κk2oY0��镃wr-Hu���gMi�Ԡ3��k|ݔ4Ў!Π�����:�)�(|��X#1��,�"9���%3}�vv��f�H��!�C*v*�t
��������Z��M��mI�G�~Ҏ�n��&���#ۧW�).#WQqc�K�7=�u�يԟ,�v%�T[wD������&���&G�H%��ꈤX��2����I�	_��D�ҵ�y!��qU����(�8D��p���wP�G��z��!�$��S�]a)�"R#M��D� �L4{]$�h�����Z}�̄W��Ѯg@�|��[�pj��3�O:�bvxzR2U��:���]��:-b�L�]P�1�W	���9�2��VWQV��)ǫR������\�Z[P@PW����a��X"�D�V�4�m+���E���y��n����S����*h�s��SA�!��H��L�=��Y;U�sydgɾY2a�쨍�aq�(.�Vx���ň���t�	����.<�i��h����	@J�N�.Zl`�|���HG}��~�v����Ww�i'�x]m�q�?�a�AU�Ce`����ϋ��jH`I;�����f��� ��Qu�9E����h|�bAְH���,��Vg0���������w/��Jkp�څ�T��~=`}�EG�6⠭��Z9�f�G�	�㴹����Z��N��8��-.^� 4�Y� j�9��[�0\è��\en]*O/���R�Q�>w��sA.A��"=�i�w��C��7�)����7 �W���� Ӡ�s]��\�hmV0�z�3A��[{Q䒂sya��:���nhM�$��%7�����7�J�� �Oq��7����-��S ���l��m�)5r"ߌ������Ӯx��u���	����9T+X��c��6��y9yK����h��o�	9��w�'|W�;bP�|��%D�5��]����3�j�z�_�ߘ;]�����J. (�Ju��Ap�V������>i�۱ԙ�vYLNF����¶���]�����ǒ���<�������ζ�H����t:��Ҵ7��k��	�2XZ~u�Mr��S���{Ϻe��Y/�m�c��S�hR�\�����XP/�k7/�����@���3�V����g��z+&#.`o�Fݷ,�����1-�4S���b$!�ޖY���7��vƢ��C�W^��!Q|M-ˆ�~��*�2o�}�� A�c����ߨ�?�_|o�.��y���J���$ϘԻz}�b�]�K�
*���;��{H����dj�ϚO�ćm��+�*4�菃�.ZjR1X�P���p
�CB�b >̙�E��>�Es/\�<&�Ou���?[�u�h���f,��t?���Fl��h�@��W��I�����~G�J�� �Ѯ���yKٯy�BFg*�$ƅ
�����}��FἩul���(��S�.U�C���P_�#Q��x>�]/S����-�=Ӱa:�@�7+��Rm��[��@��6Owx��"J��|�K8�: 7��ϙj�TDN1�^ST�����u�`4vC��]���pq~@̶�AYk�X�9*�;�����u�;]���)��i�#>*����� ��_���#���å�R��1�ᐲG���B��5O)`[;�t2�.��[�?���ݛ�C���i�j5��S�����J�GU%�j]�<�HzdxHn�vp��Ey��E�H��կ��CO�����������	>/��� ��7�ܐ��HK�4<�-e\���U ��M�����KJ���mT�B6�t�S�ĸ����$�a��Q$\
��q��8h&1qF!���e}q�)��(\��}��'�T����O�~����)̯�����Ww�[`�;�V���q�pS2�����ذ1 1�??�E�6h��YA�@�/�H8�	�ė�=�k��k�V�j۫ɜ�1�U�3�O���ä}{��}�5t����W#ض5�J  ���&��$�p/�9��:ԇ��p���H��+G�vo�n	zs�e�x�1[!j9�:�^J���Os�1)OYp��)sT����b�M�m�J����aqe�LB�YN�;�X�:i�}�b���I�O�$9t��:�@�T�c� z�����ubp!�K��J]���נO���pn��'{�hc�-�]�|_=�7�5Z��,�zӗ�=�8�����΂Rԟ��������
gT��:؇��	���Y5��^
"b����pA~�b�p�1�?�H-�t?�d���ՠL�#ۙ�<�
,y*�?J�A�&��p�r�����HhG��I���Rz2���[��5���Øv���j�M�xKfr#��l�NL�(����Ђ ���~�z���w�P+^l�DL�MSbeb����%vqQr�"���~��9R�F��K����?�f�ⲏd%� ��ڞ��_��mi��}+oZf�Ŵz�M��0Z/.{�}.���i[������F�%�˝�O�(Xr���K���9��K��m��#T�ꭸ�W歪f�� c�z�1�UgIoMn��r��orx1��j�ݺJY<�x��K�?��))G�Yd"&��Ԛ@ަ�Z�pc����W)�f�p��_������^�ªB,VB��L}��	����75�3���ڄx��Z��O�O��U���Nc%�C���6�ŧ�CI)5_,�x˧gH�b~w#]��z���Rf�q�b�Dsw�{я����R�6O��$��X����:7&s��%<`����ݩ�Ǟ�9�f���"h��q��3�אh6��=�5p�5;�I����W���=�?��������ԅS2��;�p{�y���J��X�iZ�<J�}�YΓ�$�d��'��\��@�sS��S��3q[$�*Ǌ�'�,@R�~���~�i��E5�*7u��=���������G*���h��5��R���>�5��a���f�y��G�}CK�~�Y����{X��Z�H� ���H��˼�F.^��\^1v�?����t��_��n�T���C�H�'�}�