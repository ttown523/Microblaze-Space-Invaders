XlxV64EB    fa00    2eb0E�'3�l]�
C��i�>��h��6G"Ś��5ۮ��D��4�[
�h��V�k�<0�cR��\!J��+��FH��,G�_ ����XffP�-��%B�����KH���X������ ߴ$�!�g�A���gG\-�8ݍ�8��Ҥg1<��#p������M՜@˅�F"oQ��fdTpE
[~~͙0��V]WP��vn$���lٚ�n(�����ȫ�1�Uc�;��Ǩ\Moqh�8�I[�Y�v�D��1ī��7�ˊbVFE�DR����-`�ϼ_ht�;����a���%�.�I�.�����O�[GQi͜��Q��(m}���HȰ(��u��<d�sz�o틋(QO�
:d��������U���M��HF@j�����-=#���x��;���~�Y����櫧䛹�u%e=�B�Y�wf}Ķ��{v�d��c�׍�TA&��[�FZ�Jn�E�l��`,=�+��@�s��(8��l�q��ն���n����ͮ�S{��~4�ՈzF E����i��v�i���*�Sʧ��a>_��h���?,��GШ]a���_ÐY��3�i�R�f-�.u/E�R9=)iR'�kԧ���l�[�5���U�3hLA�?;��Q�=�Fmv���GN`9�ziO�?_����Ο`�q-�[���n���"|�S3�c� � �h��ST?��,R�(k�8��f�㴯�+=a
k7|F���q�QG�8��."��>��^'����o�;��_��D=@�mTߥ���U�!�^g@1/�\Ն_f}D�e�s@�I��S�l� 9��_@�����j�PkT�� �Ҫ�׺�(' ���k�R�n̕�ٜHX6������W�x
���{�N^>�#G��C�^7���M��mg]接s����L�;�<���D�]ɻhs&���[aݩ����=��W7Ǻ{���pc��¸�Y�����g5��U��X�� ��;�=���s�ޮӊ��`g�='pŊ����p}����!FI�̙ry��{�m�^Abs�?�kD������h�I�j���$X�S���6<�LX*�O��	M���':��Qq��.S�Ku���v��J7F�W�_|3����p�Q��A��H�Ys�e�`M�]�A�s2+��`}�Bc�������DF�^p�p�/)���$ J�l����+�Ź3��<5�79W��I��J�(��:p�� 6��#�q���DTI�� �Xh�l2�:�h,���~r��D���O�*tr���1j�A��
�6���r��M�oQ��떎pT8�ER�yz��VD.1�8	���ɡ�FE)�'���@i_q5U��ܖ�Y?{�~˲��+u6Y��f3���{�'M��H����}�X]d�����}TK�;���|Ku;wg:,���NCR}H�$��^'��Dq�s��`��-
*���j����1I�\~ƦsR���jJ���w��e`��ݡ�f�D<���� �ɠ}f���q�ND�Y8���x��ϩ�&ߤzT�!�[j�Х���R�Fu1H��5��o�!Z�D�r�
�s����N�e���cE	/�%�+���R��4�g>{�ڊ ��Q���m��/��Mh��G��I���߿�=�J����t/���%�f�&`7C��8tjz�EK'g��r�n�c[�X�7D�T> u�P��7��s��һ��K�C˼%ą~�#���d��,�U�H=�����|��=�@�_2�O�����x��ۺV��&��/�H����t�m��])��7�#�ۨ\wYz��0j�y����`Ő�hƵsN���>�G|2���vD�"
���m:5?4~�\�R*�ĺH����|�_F�5-ѻ)�s�х�i�����:�
�K$�?ܺ�ͥ�TK(��*�<<m9G)�/��̕l��P�l�G0b�*�����"�t���)��S��VΊ>��m�W���~�[&���`>̎��������(�(��2{���W�^�$@5���L0�< }� T���0)���(z�J����sQ�@!���|Wtw�R�Ah	�Vj�����^t���O�����)q�)�Jl�U#���ѣ�Dڔ�m��!S����Ƚ:���$���CQרG++�|�h��	�W�-�{����D���'��	��"o�Z6��S�v\c� ?;�_K,�f���L�Ԏ|���]u7]F���c��T(�eWAJ5θ�D�"��%�{/(A�&����8ϕ�.�1�jm�
��}����ս�6�� ��f��d�֊}%����w�[P���<�2�[c�?�[x:�͕���^'P$�:B[}�+(.���6	;���x��p'�����GQ^R��/���\�� v.;��g9,�:��~�A,��(�'�h��g��zkkL����=]^�7s
b;��*+�=F��uQ�-/IG��CM-��@�0��[G&�-��A�'����Y�o��1X��Ք��sL	<@%'[)�5��z��RR��a��.�Kz�������ք����������g�����Dv,�=!"��#�!�K���,sW�R
b��h������.^��üL�WK�Z����S�G7E��$�7��ʼ�W�L��$B%w�T� 1����</�������jO�}�]��I��8҉�3�`��u���y(�0F��\��#�3�k�T�υ��ʫ1f17�!�wh3P/�����Q���_�!�w���2�3���վj� ��r9kqF�T�q�eb[�z�И.���<we������&}�k{AZ$�X�_�2A��S+A޹�j�S��v�yb��(։us�`h=~��\?e�?�i�v���Xc؀�����ʏo3�84dh;�G�M�� 8#���x��r7V����U��h�a:1(���]/		J�7�Kp�k�B
9�&���q=���J4~�c�W�h�ݺ��y�ޏ/v����L�x$���{[V�ض���L�D�%� ;��B��~��O���p�yގC�H��ցTo]�ϕ�����4�Jx|����B�;��zwS�mϊCa@���Ё���m]�)�6�8�v��1l�HX֭�k[A��9�W�$���xP�8H6R�+�ӧ��l��LQ��r�v�,04���Rd���'�C�Eq�q�6�9����Ĭ��|Gd��!s*$�@��/Ǚ�^_��@S�G�q�֢}V��2�5j/oZ�=a	ۍY��9rS���q��?��ǮY*�ʦ�����ZG?57p��X�ն�ښ���=;/�Ͱ�tO��kT��t��,������W?�Ѱl��gÕ�����VF�h}��gv,��I�(т��ѡ�mXW^��$.Fn2~��=1n��jx9�w���^��ae�J.�`s��O� �6H`,��i�| E��^X��KL��@ɬܒ�2*�&���>�A�����_�w띧��v�g�вl\�Cmy4hkуF���0+ί�E��}��F�`��s_qI�|v�u�}�j}��*�.�WAx�j�6�5B��b�-e�0�I�q%?^&�@�vg�z���g���aU�W�������ϵ{+#���H���j��W3��Ō��/:͇��O�7��M�B�d3����)��"L��^��F}|�#Il>�ˠ1�sb���&��Q����ַ�]z1\+=`阯.�6	����d��-5I!���)"�.ȣ���@�_	IS�!Ũ�|ܫ�����"�p����J^q��j7��uqc����oi3Ɓ��p�ҝ��a��*]hƑO3d��^�5�i�h���f��/��=Ǳ6����^p�����t]�W���v	%��C[�5�v	G�
,���n�W=ö��	�N�g�)����]m���p�ʋ}�ě�/��j�Mח��/*�&�]Ttb���uԪ-��fX��0�Q|��p����	�XSÝ�"QtVE�� z�(	�N�熡ɐ���ʞO`m�u�v�B��+�g�����&�Fh���l����g`rF����_x��ў�b.W�+��c��zg����Q,�rӰ�9�r^-+���P�7���G�#<p@`H������}�,�@�X��*��YLy���f�B
@��g�1�����.�W1�Y��.f�`wX�>2l@��m�[�������#t�|+�tک+�*J�b�'$Ɉ�$���s����a/$�ЖW@8��낧���K0��R��48�]�{��ޫ si��W,�\�;�Y\oS��yBe#��:�o��H�4�X�d�r8Z�zA<�vO�aP��n&��$8>&�4&h�dJ����Z�Re��S6'�-�ᙜ`�� l�Q������Z����nunH�s�Lz�Գ��!=K�2kp�k�)"Ie��	���-[!t�=0���F�8jl������Pe�nn»JB�Pl��;b���_����5Y����VeM���Z��}�8	�g�Y�ɺ4;��$�I���������'�h�I�ō�	;�"O��M*����M����I(".+#��� q�"�<x��:�� ��I`)��lp�΂����^��4@3-$Ԁ��?23�^�הߌ�&yhB݌��� �7WP`x����5����a� n`c)NQ.C��t����l��\����OW*���f�n���ƴ2��(>*R(�T��r<,�1��+�	���҇i���>	�~���ڮ�D�L�����w"'Q���{@�ZI���{?���UM���d���!0���0�	S~j��Zm*j�՝�#��Ǉ"Ļs/|eQeBޚx��1S�ňBb,i��l�D����_X,�]776/�a��`�?��;㸟ܩ���5�]�"�ߠG4C�o�jG�O|�*2�L.�sa�ɞ������'Ode�b�?p��f����vt}�v�6��|�r�%���}+-��X�kPt1�PI��U+l��W�e��"��:�K�h��)�f:<"��G
��f�S�+�,݇��=xi�a�2FA�!7�ԇ\�k�=M�h;0�G���N�[��-!H���3�\��b�!ngQ?O�®�l�Eǲ�pB ����F?� 8��'E��?T����A��4	9$�H�c���g:6�h0H��/�qx`f��Q<��%UTp@�4���jKS������5�����>�ۅ@�h�������]<U,����2
��x�7����r2�-�N��P�?J���̥D��>�+j~wZ���"B�>DJ;��C��7z��l_��$������}1�_)g,���B�%d����/PJ�e�m����~
s�\���g!&j�9T��Օ���W�xɍě�N+R�g<�V8"S��" ��3�H}�L�4�rI�.�]?,��c��d����1Ĕ���+�l��Phg?����W!��/���;��2Y�l2=(�K�������8~�Hw#�}�-��&;�P�F�;�i��6�S~�CWF�'Bbb�� �lД|�b%h� (�]�._2UJI0,�hIpCߕ��iIv��2󞠂��S�fbJ$ĥQ$z�<^gn_�m��R�H�b�C�A�C��dc{%Ҽ���;�?�<�r�N�܄s\����hGĻ=��mE����
>�q2� ��T���r�xv40� ���Y0�zo+�ǲ_��h��y%U�җ�#'�j/����a�(0\�h�ڌ�/I\���>
	b�7��<�������^Sl!�+��%10�b��ن�jZ�%+Y��rd��AE���	n�'�W��������PJ��4�;���ŭ�!f0�ݛ��8\��l~��5��W��ט��xX96 q��飼�w�bH:���Ng���\^��R3y�%)���Tj,��t$�.$~SĿ֚�["�¸�p]c\$�}D���OlS�1����c���/�-.����GܨA����[p!�~C��F��6��ۑ��ES�.|�PL����Ha�h�B\�kY�K�-����X*Ar��P&Q�1sb��}���Qg ��`?4�������`'uܨ\ Xũpt����3�k��A$ssy��w
*��bs�I*:k,j@qK��F�˪$����&�\s�st����f�n�]�Y.c�+�7tל`گEz����N�7���q���w��#���H����Z�W�����]h��7��v;A�8�oD^��J�p�(�0�:NO�di�$\����q��nc��?9��*@ě~�W���

��2N""���?�QH���ڣ����|�j��"���N�vH����-U�^�<OX�	��C��9;��*j�/���o����?�i�! /\�n7�f�v�#D���k�	�]�
�.�!�\���0x�y�hL�8���3���G3uq3�!���9줄������l1���n;wg�ÄV��|��PDI��fP1�E,�M�����B���p��s�R(�-�9�vq�[�2OM<'ʮ�Aw���ľ�e�A�p�S)\����R��3�9��\�%IݿC��U�R���0��&�p_���p���e`�W�����i0K�|5^Ź���}�H}kFQ�k��d˚K�x	fh>�ޘ(���\�B&�=ܴ+��ӧ�/����HX��\���+}(�$o"F�x�IG��F2���,6�T�s�Vs�mR���h�%,�@S�v\��䬱��F���t������=���،�N��6@m)z�9$�;�M�eK%�b��.��N����;�����$0��[�-�����|��9�WC�ިYG����MTx�9�*w�!�èJM'8���硔~$��y�w����@M�c�q�]T��J�i/���?e���-��|�~͢,�O�1�7?�x/�c��h���i�1�]�k�<m���o7�����n�(�i�^'L��O�J�D�K*��G"��/n�59�:�����;��m'��"��xJ�����2���˯#���m���:lb��hk�g�̇6=�"��ވ�E��Ln�^�P�� ��-�z\X����%�B�a�'�xIe#G��=�e�u�I0��tN�8ܞHBV��|�1<�&]M����,�������4�3Yt�Qp��:���J�n2�Y⇑�w�����~���cC^���~�wLUr��B��.��?H�q��T:ۣ{��{�зض1����Iı�ƬƼhnM�֙�;,J!�ߔ��3�SN��͖Q���*��:�kd���,m��U٠�|n)#�b�m����LU�_�+��[�u�t�k�d�~>�`mH!Щ�	�Dy���tӠEi��k��+��U�x<\R�
�V�T�A(��g�;)� �R�A�s��g7�qHB{^=�Y�&�����:�'9������1��QGQ�v��o�5C[��ҳ(@sS	�."*J'v⥆2����)r�'�P�®�)�˪y\���(�$�~Xڨ9Vk���?u�����?�C�R,,S =�DN�y�GUe���v�iߜޙ1{����r�U�p����`w�bHZ8��(��k�.�ڍ���ɑ%���9��B"� �b�j$�؛+-@����>"[V-�E���C0�Fޮ���`)ʈ�=u�YQK�L�n~�8��)�������Rc�g�jJ�u��{�o�5��pl7H�!��v �p��t�o�0"5��a�\�`�-^Y���"&� ���$+���k<+�Z�4D��d���eE�(& �1��Ot��F���̖��20�ς��R�F���f�zPq�=�=��3�U��MOt�o+5$���Ǹ��+7�X�5Ag4�ԿWv܈,�:&ME�Ri�)�Ǥ��Z[��[F�^{��|���Mm0�e��3Yncw�%{��Mh�u�c'.��t��}8ŗ��н�ʜ��?�i���G�j��%1-�M��	M0da4ʑ���Ad�G�m\�߬������ǳ���-&GD��RU�̵̓�uC?vD�[�o�����E��˺tw��<���J��DjM<�1)�9�s�wPS��sD�hT'"I?�O�b�
�BeݖGWmP�6�������m�Qm{�
W̘�߾��,�_ۛ���*BG���2n߂��_������l��j�z���ȇ�<���{<���	uτ�E����ST�+�S; X;M�����H�^%�j���!�۫�gX�LWw� � ������e6� *���Q�&%�6�����vv�+�Dd�L�ڔ�D��
��M�y,Oe��Mv��
�%��U�_��>������]Q0�Ko���t��
-�O՞�!#����~����Q����ڻ{��u���|Ur�H����?#QF'�Q�E��U�S��I(�(��A��� Bd�a�n�M�c��n>s80�h�t�Lab�imb��ɱU£` ��7��J��Z�ݜ��=l�(��H����	xI�Zg5��?#ȋ����K��|��	=W>��D�唣0�5!����KE6�
wP���M7�u�P���?^U��� Z�{:�a����\a��z�W{�[ڻ	�4��2�k��8
��y��v�_�Կ����]r4��\���V�Х:=�r����[Pi9� �
㌄���^<��إ�s��R�rk�%N�Y����:���$�\ގau�p����J<q��514�Bj���/u�;����e�\��@nk�8��a�b2X�����Ky�s]�&8~/��kg���	2F=�'<�N6����!�}'�PJ��� W���	�7J��F�VÒ����A-�=Rܟ����`cx��:���Qxs� n���l�p=��i��=C];�<e7N�����|��o�[�h�
���eRb<o��v;�am���Y�H�LԮ�~�[$��U�̸�����`ڀr^��Y��-���;��힁mܢU�/��	FL���-��/�Y���zT��ū�5*<���M5�<(T�F��GUB�M��#ݐ����-<�o��l���P�9L��� ��AsQ�Y�I6%�%��x 9g�z8�>��dƅW��A� �!�9�f�R���n
��Ҿ$�?��M�׈Ii3/���=��r�:��K^Q;\z�[%`�*È�(a����zNwvlׄxN9��H`ao��'͜�	���}���Z_o�q0������g�C�����\�~!��}=��#��\����$����rz�Ҏ_U���(���hƞ�ˆ����m��]�52X�;�2�yZ�H#O��IC@F��S!��$
�1z��<��{-�B�u��mb�C".�3�1s�n�M��P�ؼ�	Ū
�RJ��WdPp���A��M�N�i�d}'	[�?0� 0�����2J���k�2c���;U�ZiNI�6Y�/.�/��>��A�oߐhE�E���(: 4����%Lc���e04P2�~�/�tzk�@�̔㱴r#n�Ah	�}����3�M�d;���$�̄�I��u�q# WjR���J�W3�**O�� �K�L+??��9���/\�����(��|@��2p|��5Rw�J�2�l �����ϡ����}Fq_B�s�O�6�&ߘK�9P�~d"�e�`f[-������z2ǒ�ʛI����O��E	a�YE�����?rE�D�ΖO������>y��˲}�<?U뫾b�^>a�3%�4�4�FLEߒ���@���/���G�%0f�b����Δ�����/	�ѯؾ�Q�w"B��R�&��M&J��г��0��̿0��UGf�w�i��D@�$�.ϗ4-x;�
G����j�1d�F|��P��9Ĕ����sk�3��潴����ɨ�����n�������Q���Y��!p"���Ueo����S�zn��K��L�#�����4-�&���@��k���|��~MDh|Ea�1����mv�"���!��	d����B����G4oI �����T^�\�<��g�2t.$�%h'���g�h�������&�_-:�����Wy�N�v450E�3k�e�|�s�c��.y��H�YO���}�G�<�A��g׭�\~�\f�Et���UN��j�Em�+*�V�E:/�oZ`�t�RퟛN<8���s�oa�k<GKFgx�-w[|ʕ��ȘG@�m�g?�����	21���,XیI�ʛ�a���,���Ɲ���6�^��� �˃�?�vE��c�\�����頳��nus"�~KU1o��\�Y% �A�I���+���{�;j~2k*�����#BI{DlI����,=��p�5��;5���BrM�|%�>>���F�=Z@�C�����к
s�Eۅz���k�� �Ɉ�'�X%}˃@�8�j�N� �C��KA�wқo���/�ȵ+rB��ę��0����2�A�5t/�y��LC"�$��\"Uw��0غ��4��c��&ԣ$���	v�7r�+o0��vX�A{U�Ӈ��CX��:�i��$��k$� �1�$(��8��B�\ �]��sv��:�W|�k;I1������ ����o���b2hF�v� �_z�*T��{�(ʛ*%H ��9v�1i2���XZ� �w���Ɍ�R��zq
b�J1V�������'�6mBuhվ7��-�3�i1���7F.���*�kev��K��N9/�O}N�߶z�������b�����o3i����4���6�n�W[�Q�G&^�<�n>^oÞ��7�$���R����a����7?�?��	���Q����J���-X�)5�����x����*��)-�7���['U��(�� ~I�^Gr�J�Dx\��]���Pq��F��Az(�Q����x|Ҭ�����H��ʛK?�<y3N��I�S�@u�	�tI���b�Z��Y�+���F1��4��`Rz��b�>L_L�H�H���[�e��(غ��~p�8<��I�er�#�Ƃ�J�e�?��jw��js1��-�_�La�Fr��q�O0\w*��W����Z�������g���xOX���XW�bp�������L�s/� �L��%B]!9�{]�N���'�|<�x���zy�S�F�1H�]8�ԥ����_�J�p�ܯ�2��[��u��HS��Q�gt�0v����LjS��pc"�b���, -N�#D�nps �����:�"�%�ݔ�%'��շ�7�/� ���b��p�&7�gfIk{��O��2������F��1�.n�d��g����'�ʶ���u/@�v]�f_���	q�dc�Jr�&�H[*�3��7�G���٘ƳĶ?�cl�0�]2b��C�ҕ���8���?T>LJ�i�0�$&���CI�����JLx�vZ�Ǖ���v�&�W�Yߕ-Y��$Z���:b���,�G�:�a$�Dg��m�\ɪ�Ť��`�ꅰH����.��đ� �F�i�Bdğ��d�t�q咤0ɾq�}��!T���C5���F�X�+& '�A4h썜���bd`:�D��JЁ1��>�vt#k��q�78�.�v�&A�E�:�4,+��7�V$Q�^P�� Z20�L���?�΂o�!A�-#@~(i�gdK���̠茟��yM3�%rX�~��[v���&$H�"����͍�^�B�&���Hl� ��:�<��]��s����>.1��>�<P�:2����B���/��B�E��ߪ2��^���3p>�^.n��S��l���ܗ=QkH�p���VXlxV64EB    fa00    2bc0�g�H��9���'!}�0�w4��9u�[�)�����h.5>8]���aݗ "|�H�k^A��������$�"����ʿ���?�#a����?!hcN� 8X���c<#v�Hb�g�\'iŃ�Uo[2�Z�O��mK�N��N����(q˪��W����^޸e�?B�j�ANv ��$/>aW���z�c�8���;�v��3��n�w3D� "�2��-h]J>_d��u� r�M~;"`�䴔P�!5��ðŵw��j1� �Ið�J �A�&� 4���t�Au!3?V�y���`>f�/��*d`�P��m�3�< �se�,��֒�$�F�� $z��/3�C�Ks�Y\$NQ݃�q*�&���;�!�ɓ�H��u�e�vQ���堰-"㦈�1�e["�����K6��-��&� �vp+��"(24��;���k��s�ƚ�%��4�?1��BV�i����p��	���_�S�%a�h07V$���ci�b�R,&�q��s����PJK29<���Qx�<�� �;IX��(���|���GH���MK�P�Ecr�A�ۊ{���z1/G��H3%d����Q��ʹ	���7'��aH��%6)pT��9.���{Ë���'�~��$��jy�UE�;��$B���y�0TD�������?P��gĦ�D��"w�I�Á�F�CVr�zI�9�zӕ()t�%(V���䘴��q�b��b>����WȂi/���WX�Х"��K�^[>qƈ�u��%�ˋ����2�]۝��MT �X�A�zs�8?e�+�#��]�RN�
������K}wS��o<��r�5����ʜ�W2�)=��>z'_;����bA��䇝գƛ7}�̹q��w"�ڣ:�Ͷ���
�6E3�=@f���]ˎ�eF��̶
~?�:�r ���4��l������w�0σswT(C<�G�%�1*�;�M&q/�g�q&�x|f��h:02�Y�T)�H��	0��ކ �����^"�p���l�$��J���S�� +��f�օܦR.C�&ݯ���jrb�����=�k��?�cJ��M�k�	���@j�)��i�=�wOk/a"^.�f� \����r{�ܧc��S�ӈ^Z�-l��8�3.m�0���x5����BӔ���d��S�X�x&��4��"�h���	����~rק���IQ�Mnq�{Ȭ��L2�m��Z����۩\7�ĳ$�lBk���g��+�[����y	n��������,Q����֙��M���q�τ���>5��gV@�]V����e��hn��h{p1�ˆ����~A�9�3R���"����YBX:ߍ4Z1�c�J@۔����ʛ�ɐ�Ť�d��hl�*�cC��������8;�>S�]�1����K����?�zQ�?��L�,0����Yn�I����T���Rl�g=��PsL0��	"�m��1^��B��}��:��n2���oh)�O9%���VYD?|#��lD��x��2]�T ̲���!-蘢'�M����/2~6<2��Y��Ƴ�ե�25�&u'J�5@Cʻ	1h �|�Ѝ�y��pe|�E�+�Z�j��"���z1Z!�T���c@��1���bi�+� U�aa'�@����Z�q�!��ʦ�I��-Œh�=�J^<� 9��J���e���0����L��m��u�GՄ��g���lgc����g^���pޫ�_ah�0������.������l1Ho��I�"��':��T������_}�x������ȕ�P�0�u"2���6��T3��дɬŧ4�ۈ��u����G���r�g�H��?��2T�1D��Њ���:���'g�S!���d�d*l�|�����I��Z8z��qz�l1{��%�#"9#�	�$�Ǻl�s���x���.>!h��u�CF{eP������])s"���s�2�.
D�$X#އ�Q���)~(E*�l��k�n}�Y^��~�N]����_>��v��6�x,D�<���hg���i��h`R������e_�>��d5=�����Iʻ�4�=�It0u�Ja��������$L�-&�+�7�����M���V�)����}�$F�F.���<rF؀.RB�E� ���ӂAU�\�r ���+k}��I8���lyZ	P�)�pI�[3�P:Z��t5�ַ��r6T�x�6O7
��'ގ�Oz/N���Fa�e��߰���V�5�y� ��<*9���菾�0�9!��bK�6OA����b���4q�O�?&�ef�<���mO	��[�#�S}5R/$ܳ�W"#I���+ۜ��V�X��q�<����
U�Ǯb����x�AM���՝+.�X|�/ȵ��s-�9���J������fK�n�{Ʈ����$@�W������ԋ�wzs�����$,k��#�B�����!4}��%�A���ᇱ+���p��>�M�Rʆ*�J@j�p��ˀ("��C0����5mr��7�:|��'R<����y��jSߎ�S烽��3�	P�od����/�z�d���o ��)s�eZ������}����?�T�=W�zߡ�@+b��m�"0���;fh�d']�=��4��f��A5��Jx�0C$g�y�6b�JP�F���n#���k%ea�e{~M7�ꇈ�=̻R�7�_�4T8>,��/�5���GX�4���w7���t���M3�x(�z�,�_�'8��bH��';u6љ7K* ���b���pycf#9UD���f��nJ���|�EA��o)�oBnp�k���|�س�;�Q��@��x�t�v�y���	��Z�K�zR4$�u�d58�������2�����;,��c����a���ew�}�� |��ڦ�͡�1���=!�%8��K+;js��P�F�y�� ��,�H�:�&�u�k���o=���?�Fo3���ۼw+��|[�>UTX��~mу�/Ԝ*����4�w�J�q#���!���nA+,���]��8ǌ/�,zוt�wz3y���;�K��wB�-�-+T?S�����
��(}:��N�8��\�t�f��ᯅQ��p���F`4�����u�b�2M�W�-+�f��ѷB,��k�˄����*�
��������H>����!1_�G>M���-;��4�Gd�:=��S��6%�w��|H��*���������}������p��8w�����c���,ե�l�B͉�V�Y��	��5�I��#o��K�z2�����
:����C�y˰���RJ�A�M ���:ETf�/��M�@�:T��#��`�H��
����(۞����݋H���iu�|��I�^�}�@���V��*Z�B�_���sbH!$~6�B����6uL�;ر�`iHE�"2`�xܼ b��]$Z�sJm��{�����L���8�&k@��";v6��-	�~aSJ��L�t�����ıf+Vs��1�r���|���m!.�h�d��>�/��j���fP�/ŕDR�CqmR�(ϖB��E�uzD��ws-���YGi�
5^N
�q1�5%�;�������h�(ϣG�-l]5N*2s��K�<��9Y�No[��O��lOK$	�{z?��9=�ϓ���|*��n-ap�K�uٽɼ�������P;�&f�<z'G�l6�8�"���p���om\Kr�4۔5\?E�ʷ�6c��q�i9��ژE֔Pt�8�����9�I�D�G�-9kb�������^����OzI�!Ԝɜ!0wr�n;XT���.M�R?�ݔԪFá��'��ͫI�zp��f=��G�G��ka�S�{'��*&'g�A��
�]���OX�+����bF_�2�c�P�1*�&�%@�.2�O�щ����k��P��: _�"�lԓn�>!	])[��t�i*�2�f��G����AV^U���Q�w ~�	����\��C%;W��!��A��Ʉ�웽Mf�i֭$��@oq���[-d�/��o؅G׫��	��f���'|/�����������T���R�x|ؔ�m�wS�%}�y�~�C�]�����!f�I���Q�h�u�2�x� <`sP�3_��*�t�A�ͦ�0���6yQ3:& ��fl���+�7�z�>�
�t)����'��?)E ��$�2�!�Rxu�I*�0 |�K�g����r�R�
w���6^j:�jU�b�0@�($1SͿ�2��ğ��qrzy�k��:�S�!�c����%�Q���-��z���G�}�(ޕq����������Rx��uf�8��q��U��n0$��6#�I��-+��K_y5�v$|gp~�F�uK�UB�į�za̘�|�ƬG����ה.����B�6�.�H���e���3m�G��&�墆q+W.������( ��c�L��*�IñMX��@P:K�p�(]�*ꑔ,˼��OU������>n��J��^�/^<������:�]��7��4��i�h�r�R�c�͞�!u"���~��U_O�����!��X�|ؒE�͠�ߓw��Ag̨8��w���bS}I�"-���/_eh19k`��B�?�v(q����6����Ո+r�	G��Cu�9�A@��/u�P�����s�V�ʟ��$864�Rv�e�.�fW�Qޒ>�&9��U��N���0k��I�|M4��ݛ��ݾE�LQ�7�����b����&����B�gg쬐�R�%pW��e�<^�
�k���?6�J������9[R�\&�D���U�S��
�S�L���>��T�m�����O��r� ?�b}��?�+&qx��ƩZ�D��Zg���|+�Ri�((wv�c�(�JZp#ֽH`+��0n
&�B��^���jIh;�_e�Dǖ�b��;��8�;��ʩZ��n�{��)9H��4
O �6��O,�䍮�i�SǰYd�� s��#��3���D�>��S�ܳ ��H��\��:5�������h ퟉��˦�Jq�=sI��
&�,��V�ڪfHB��̧>���Q�Dޠ�F����&t:�d��s���I 3nr����8�ө��Dp��0N� �\h�hy㆜[�NJ$Q��Q�x�	���H�63�1�� @�T�-�l���ˈL�&f�"�_��u�@ x��p-������N_x��1�)�L���R}�ḻS�zW�[g�^FZҬ )z�5�v���^�
�ҡ$�5i�v�63�Ԍ�jb�fD�`8�7��XJ��O�wK��#��(!z�$��W�w��y��{G�j�K2[��"ZGKna���]+pj���V8��n��z�qK�^�ވ��}����)�2�ػ�eN9�� �F���:�G��Sz�����k�������'���� BÏ��}�(��
Ρ��q ��E���L�
���1��\��l?Rheס+:�����c"0���H�t���#o�)�����b$���Upe���z��A����C9����~R¸ l�!�^E����ѐ������z�qd$%�P���'`�U�jn���:D=g80��}�08���|>���.��|M�5������1k(#!�Goŉ�8<�c�PHqN�fy:�Юy�'y=�C8$����t���a����e�1��C�������rZ(�S���աN4e�q_�9T@5<
yk�G銭j%�:[`��[����6}���L��]����G��Q�����Y��ص�����.�|*�`)C������$f�NZ��P��9�u�5��V/Mg��]���ˤ"�Lj�wF�ּ��>�-��U�iF�1*�6c������@���W�A6��K���׏}ax| �V�m�+|*�~Rr���c�ΰQ�Y�_���lf�甂���g�ICy�`J*�~/M]i�lՉ>eҏj��r�*UqA���"��"]��9�PL	��z�p\�aj��62��6�� �	qh����_F�n[C׬��b����`�4b������n�f鿽�����|�n�g
?��WW�$l��v���!X�����E[��1�'������A�:NSU/�tu�7Ag��$�j	]��|���D�� s���$?I��^����"���g-zX���|�6֨�Ѭ�z	�3�d��/�Oi�u��
k4ܐ7��ZM��K
�u�	�����9�Kq���c�_��{y�2��^oޯ-����Q��O��z��X9׏�����ʚD<�w��"���ҩ��si'�B1�dn������[�h�]��$���q�@�L�r���.�O�'U�;�G~�2�Gؙ��-�#Ձ(����H�Ы���M������#_��|����4V��r w�f�q^8��hV��Xj�ej#7����~5�}b��Ϭ��[��t�����+��B1��[vX�&;�JE&�υ�Z�|�LkM>2 �,�,����C8��B��`�#��KUvݜ1Uj�;�_�]`ζi���~��-q2�����@����T9�̙��}a��x.�\8�a����F�y�3�蘢M4*:9@�s�9��akC��_�����v`uWU���~f���t@���z�G%����cb0�SOp��b}6���'_/��"��?}J�L�i���V��rt;�_��&1��gAU�k�z���ˑ($y���;�� �N���	�Q�5<O�#6��g� ��_nj>�ĖPO��NN��ʨ���- ��X����9�'˅ߦ~����\�7%�*���F��cݤ�����{�w�\����S�PWX �z��dgi"�K����܉ܶz׸��9� ��b�{�=w1>�1�I���g/���E����Q7�������L�QQ{)�����o�-i���(�; r�O�;q�$�������^�}ӌ�ţ�5.-��R���9���BE�e��̗�څ-#Y�i�X���Tc�Ȯ�ب�*�?(�`eh��ϕyK�ZCr<��c�-3�J��˞x���d��깻�ܹ쮺vZ`V�U��~yGQ�{�7���-{q�4&�X���
�� P�i��J�����b�`e!���Y$���W#;��ά���+1K�G��W��P��C�S�k��lu���:�=DB��VZ��Wf㌦�m��c�V:ŀQ�q} c�!L�|-�IR�=W�	椬Ҟ��Bf$���?N����Ӟԡ�
Ҹ�����Wn�}���LkP.`:{%����Z@ЀƂ�R��А�2X�=�H��4�K���NP/U�w睋��G�'�r�0i�IZ^���,P ��;� �7g�1��^��^1�=5�9�/=}��n���}�!�X�Gf_Z��6f�P�TE4-��ӂ�+Ū��79e�[N���
�hoG��}L���#M�l�ǖP�����7��� �<��K��p������{B�
����Y�O�d0�Z��ā�K('�Rz;z�Yk����|X:&>{f�ˋ��fi�z�Z7���¾��u�2�A���dțs��6��Q�$x!��� ��pwR�F����&|s#�ڊ������Z��;���v^�W���~�(�Y��[�j��hOv��خm���RY5XO/����|r�_�!t�n������R~�ɫ���; �Ӹ�n���0��|UL�`�1߇}�����X?`���"�܋0=�y�rN�W�+��*9��{A)��M:@�{P�5�}���!��E���]�t�`��g��,%�=h���ߧc*aM����O̝�����5L�����ÃnEA�Y�GRSv�	��X����'l_ӷ=��o������D5R�ąN)?���A4G��B�ܢaf���۞��4�mGӱvQ�0DvhW���ՙ���iA��4���WbRu��is�"��>'�y��΂Y��rQ��(�߀/Q�)g����&��4���H=IR��8i�PyL{tx3ꋞ(?}竟:2�ܠ���}�*.)����,�}I*�ό�g� :�?��Go�s�,~�H��t?ֺ,�,���[-��Z�YG�8�j��҄�]��m|R��g	I�C,|%�ؾ��x�#=���`�W~���pc��0%}h+%�g ��!'�6�U J_��z1�X�/O���e��<`Gw�>E��%=|��&����BZO4`>k~gE�{�x��t�(�;I��ɬ��ss�Ў`�ęJ�uj�)���8��ѭ��S߰1w�PWe8�x��H����h��
9��a���6�B�q-�z����1㼦��ş�L'��z�J��Y-�^3���)�/˲]�Om�"�4Fؐ/��s���v7=�S�[|�?җ8Á���_m _w��u������4.Qf�5���.��7ͫ6oz
(	��$к�}/]�	C��|������4�@:����}�_�Cx���2{�'�R�sS�w�6��^Ԃe���⃧q/�B�3��.&#��w��?1k�B�n��(?
8y�NAΊ���Â��n`$���������J��g�-�L�.�/�K|�,�1G�f�g�����yB}�2N����P���:��ʴ��c]�Kk��!���`���|Le;wB�]L5����%7���3%X3�FI��ೀ'��r�{�9͙e�4muf�t�u���� v��y�M� �V���?�I���xA��ßY�d<�<�ÈN��L��{|�w/ �+�,�)�uw_>�0���qua9�����`�
�B�]����2ǹmG�;G�{�,w�=B��$R�"8UQt}��eʂ�O��R�R��L�Ђ<�����b�{������TjB��X�������Qx3��5U�����d_����y���l`���`�����.:�E��l��|�M!�MV����C�D�_U� �z��!�H�2:w�A���b�H>�8�8�?p���ýV������]��EC�oI=���)�d�Q��͛�S�>���4����"��M��d`h M��;h�(`7hM�����A�rU�D"�D�(�㊙����G��f)B�mO���%�����(���-��>�%IGp��g��)�)\���c�ュǍ{\I��	b#S�/�NK
g���exWa��I��K&}d��}rx��^�ka���O>Ž����Mw��e��ky�1q ��������%j�ԕ4�Oan�/�$�X~q������yy�,�������S:b_�~+ġr'�&
���=��푾��p�!�(���qG�ҙ��E��\���
��,� c�j!�?1\���|(���w�\�v�{	mU���`�Z����yȶ�R�D�����N�OPR�W���&u
*b -�!�6�ef^�����o����>LȈ���0Ǎ�]�Ϩ;27����T�u�2�/İSd�V[e4��Re�>���O���E��K�%�\ƭ�m��~Ƚ�����b���1|�dch&�b���$���A�����dDh%�a�'Y�O?h��K�opZ�� $�ҏ/��p�����^�
� �,�$���S��]����g��ݳ]2So����؇7�����
R��|��~|0+f9�����z��~�H�ϡ����v�(�R?G/�mb�Jnt��{�A�P�_�sl���S�b��9lD3���E�1g��TD@�G5����w\C7���T���yvb��:�E�Y���c���L,��8P��B�������q�$��'H��$���֢���{�@6C�4'���/?�J�d?�j��K�p%�^��g����b{���*��3m<��x˦_N��G��˨�-hCE?$S�]x
�#`U�Ty���rC瞤_X���%�Rَ�K� ��y���I34��<�������z��I��|"O(/����0�w�.6
x&�>(�
Иڤ��/+��̴�Iì��-����o�Y�L�F7���x���CU ч�"
kr����2�#�H�1�����1/ y#���1�['"��xW�߅����z��Jf������5���jۀ��H?��5/���햡���i�(0�Y��*�T\8�Cr������ڏ[	��6Ώ��i��F���I��)t�N��E4��f�r4bT���'
�JO!�x�W"��X�������j}�g΂��h	o�7��&��Y�|��
rŀ���Y�aW_�ڠ�'�r��5奦��r#KF�WR������hz���D�o��E�}���dm�:�nA������5���]愆�Ma��H��/��k�5e8�X~
HX�K�U%0탨ɴ�ӱ&���W�qn3��振i���ϷCCz�2e�J:'����oMK����[��WL�҆Y��W�r�����:9HԓTj��`A�2/���#��(�M{6��Euprd�hg��g��X��+�TWm<��}�h��J:��0/
�j�=���|qF�T"Y�e�Š[��[������am-��� ��t9B�
Q��`�S�+1�㓇@�C�\5nW��}L�Ѓ#���W�E�e"�0��Ȏ��V�~�Q�$G�>�r��Z���>���/��DWRB'h�F���9_�;8eá����K�z^\s)��l���W�71� ���7���zMU�b���%�t�9�ү�
�$$B�M<Vҝ���������F�w֚�K�ksn��Y�99'�v���k����*XL F/!� ��(� �o���X�������U� Q&����#�ODu��j�>0�E��B��D��@V�꣦!u5[tm'�q�v�L�W�%
SY���>�}�C��l��N����J����=O���*
Ic.�<:�(�}#+���#��O?��C�i{�^�Շ�^�^��=5g���m#��l�>�J����v,>"L?M;$��en|�r���H��u�.	#}B��%%�+�zJ[+��ߣ.�%e�h��]�+tĎ)J����*_�L�XlxV64EB    abe1    1cf0ʱ׿�*a1�Ay��ƀp�Ro���> ���J��o!��i�^1��̈����ӄ�*M�d�I'4�Ş���oH�l�C�����g��e�7�<��ϛ����1�$�P��2�����+Q>��s>����0��9׺v�K �-�ӵaz�_ed�8�§���)H|���!��|m�8)��	ݠ�u�$Ba� ��Dv �zI�>��>�$�R����}������*\n�_@�l�������px��s�����)c�+d���?fް9R�����h���n����̴^�R2�Np0�f+�"��_T4��L����RL�f��'68��Lq�Ѣ�]+σ/��o��M^#O4�CjI��r�'�ۑ#h�_ɭko��Tܝ4~*��8��3�p����N�Ai�~��(��`��t?d���2��6�c�탨�L�)f�`�У:�I1�j�[�J=�����{SK�,����J2�nG�	�7)�?����vĤ�����0.����scHP2k��H�!�]/<cٗk��[��-��B��+9e�B��h�8De�i3���Ҽm�SҮj��x�+/ k8a�D�zū���2�6�M7k��� 6%���C���7 �98
�Kĩ�Q��ͳ��S�h��U�y�-9s%;T}7o��˦�����jt.���:PB���۲us3��Q�>�yhmR�n���s��@�fIa�3�t7Nv�%�>��� =���o(�}�O5�kT�74de��7a0�g[��E���Ji���r/�����A�L��ȥ�N�����+M#1F�J�:�*!�{g�s�"X+�q��z��l�f]a'_�jCEu�z����Bޱ���l�S�Fhȍx"2Ø�&b��\�P)E�!��E&Ed]L���Y�ů>/q�RX%~~���zuX����!�\"�z!�H��t[��l�T�]�ȯQ�<�w���,��p4~A��f��/��C�&�̻���*�zZqKP�n�\yvłH��+��+�!�٧H�������E
�S��6��J�������[��������uQ1�p�T�Y%�H�g ܗ�5SO��&�T�����c��[����au,�  5�N X����w�20W�!l�%8� %�,�e���e��dƀ�����b%Yb��h- �tյ�V�f�q�G�[�zR40�O{�z���'�W-��k�ߡ���!W�!��5��JN��ۥ$����32j�����v�xy��wÜ$;�� ~d[W�U�;�>�9�A�B�&?��_�	ƁU�<��%��&���f�'�YE���T�0���������+
�/Q�ܾ��]�t�P����K
�
/j�!8=^=�� ���+���S�0}��d
h,��ſ��y���#!�h�$G��~"D����=%4�֙�u����6K��W���ͼ�P��/)Y�|���n\Y���N��!�+軗��Cdw�$b�ھ*�J�,~�r��+ZGl��R^v��鑝/�qA�M]��.,q{ ?�5IU?Ɔ9̚�߇ݥN�6ks;S�~4����-|�y�zAC�d?A60}�IR)Q�4��� �yV��ɑ����Y�K/�w��}��\�./>�Xo%���k����
ɴ�6���ѡ�m`>raTs����3�˘7S��E���w(mR
\����ƺx,Op@�ŷ���Fk�Y=TжIVs|�.��br�*0y�N��4��_�kN�j3%��6VN�"ۼ샟��~$/5�I���v�P��q��=*\k�2Y�=�uu��e���A��2Q�RA�<��`[�ҁZ�U����Kߏq��B��l2h��x�����r�Xh���"۩'Aa'�]�t�T�G��@j�����KE+���?m��V�?�9�����u�k9��48�l廔.��dm��-Gr�@z��Ƴ�T�;���E�q?�;���9�P\KʰڶHC�\�M�^�#�Cj��]�T/�N�ڣA�w�4,5�J�Ǥ��KOc��I�}���mkjH��s!5|���Ϫ�!K,=*qF�/�@�}V��U��N�x:�Zb�jNz�(-�!�>(4�30<�N�BwӤ�ْ��c���>z�kĂeq��W
?;�V�������=�0Gғ���@�wu��LMN&����0/���J�����& �2E
�c�o�'�ÿ�aJ%Zt9�%w����iG��;ܞ,�iB����� ֔D_���!
?�?'(5�L7�M
�ɟ�B��J�����h3�S��Z�ʙ�F�``N�����4��i�TuRc�T�r�E\sa�4wi��r��E�D ̮�]�E]V��C�hM#�B�`�md��9��9�IDa�v�*݌��Fy�(���M�'�w��c��0g2'S�Q���I
�K$T{rQ9����б�� ��nY��;{�>��/$u b�È�c�M�-��ﴜg�����@r}���x���͍��T��[�dI�{��3Nϊ{�`��V��.��W�v;�Mg�e����#���im�}����ig�0� D��1`�0
���E�k�];��E\:�J�$k�5�q����B��	P̿�v��o{�ȃ�]��ru�r��"�"2|���ۨ��V�m��y�7qJa�g�ƪ�a#��)��At�8T �1e�I��e+trq���v���m/?aB5����w�:6�(�̃��6�V�������=��o�(5�^�����+�5�$T�o��W�a!��j�Rc��-B� �N�JZ��W3���9:�����O+I��D�^0e��� �Z]�Mv��<w����=�����|�]��]�%���:/:�B�D��jk�󀩫�#����'��Ϝ����)�K��l�q���9W>���Ƨ=ӝ�9�阎���)����Eޗ)��m��iJi���L�yj�N�Wmt0�_c7��I'�]k4��j����O�J�EM���e��yyif69q����v����?8�mj���f�#�nW�R���!ү�����O���$?t_��q	�^��r��jn��L��� X ����%�.���*��C7 Y�\�=����/�����9`��$9����˜S��3������U��i,%���׵��#��m|�:>'0�"L@��J!"��␲�?P"z0����\mΧqkVޖs�:�`����~=��?�� DBolD�h����t
�2�оR��|:&�o��ԖU��/_�U-�(�hC;���yO��6�`�	��q��K�(N� ��ahe�A�b$��u��٠h�}� ���	0�pJ�F'��oLj�Ɓd�݁l�2����I��I�f�ʩ ����r ��L4Rp����.�� 
f�e�\K�I(Ī�8w���(J(��,+��6�?׈��\���n�϶�Υ��R%	����b�4w��*���<���
�1��q�~%MS|�'O�E��@R�"�.�!������1��!����/임w���tP'Q�$ʛ(��%YݷiM��*`}~@M�$�C
���9e����A�-��a�A��%Z�A�۞��ٖ!��J��cyeR�JG�.��brk�n/X�ES��~�)�̫��k�dLdzL5Q/�KB~G��Lj�سn�vǊ�IR����k��Ϗ�$�$�^���j��V��KR2Mg�14S9î7o�m復�x9M4�O��#��.�7�����e�ef��1�����5�8fw)��� ��CɁ5�H+�I���~8�Cq[�� G�/�g�'��}gָ�D�<ڮ趮�t: $ ������IL�$���V�oiR�L(�T��sl`ͪƾ]:�3�B*SV��"n�p����w�����˃��&�1�l�!(�6P��}�pp�mfܾE�A��q���:rθ����>O�:2c���X$TW�{|�&�gf6�*j���'�iJ�>�����G![@�Bm{�M.`O���-��4�u��yp]D��z��=t�o��)�}o����ɧ�����MW|5_��ζ(��V��Hd�~�1�����!(�j�gmQ�s(D&z����@[/���F�Y0)�U�9l^��A�M����!ۢW�Ǟ���ʐ�yƲ�H1�PI�\�!b�)[��+*�*F�Z�G��RV���X��"_�R��C�!��P*��)A�+���n'CeQ�۵!��"�=�4J�MoL��H�4�.��M��&��B}�QX���#��s][س߁�(Զt�������m�C�yoc렟�:q���?ʜ2��b%����w�ۆ2�(�_��SS,I�� ϙ���}2�Q��Y����v�jSE�#[+��"����9��\a�@a���|�J�{�.����<��*����H&g�lO�D_`��E)���(u�!Z#\�P�
4�ڸ|�a:4)[4��(��e_�c25[N-Ԯ�������M�F4�������幞 iR��֍���5�R���C���eJ�j�[j�}��{n�"�L����!.��߷���T7?�=$B�&;�%b�������<-זk�������!ڟ�G���c{O#z`�k'��{G��cO~� �OB��_98�(���y�
b��)#�ʰ��!7I�(M������G|Lmʹ�=���
TjJ�����c��o�meDO�J�T�ʘ���O��0��" �~]}�#�a�z:{IB�K��;d�N�v�����zw�v�ĭ.aVgΕ��Ax��KЗ�6h@J=޳�|U�c�C��/�Y�1Z�=��z=N�����A�I~+�8o�B�-���Y1���Z��F.��u-Q?_�n�DY*j*�%@[�M�{�|��s���'\��N��K�B��&+gb/I.��)��b�^A�iMd�$������1��d����p1g�  �:8C�j<���?PwoV�l�"��W`	3�q�+�1-��P�ğ���nW�Y,�7�g��O.-�i��0���L �BYdr�^���y
�֩�GUI;�ۮKJime��s���#��'�Ih�M��FN��>T����/�akR����C�8��ǹ�0��2�����`���!)�����_�A�� w�����Xdo�#k�<.Ou���Z$�P�X�w�[#�2>�\����{���l�?���'Ŵн����d��K�_U ��zV�Gu؀�(��0{v�rU.�?�2va�ו U�o�!`�[�.���eQ��|��EJ7�v��!9?��`華��zB�T��7���֒�%Q�]�TyA�M`b�bN* �=�\��`z�?�����-_g�JYɞ�2B��ҵ����K�|n!���y�^�:��8i���Yԃ�5�FyRg����ˏ$�\+g'Wt��q�W�����:�h���,Q6:�+Ytf�i������ƴܿ��p���ɫ�����n���7�i��IW��rq�K�#;����c�o�4q��ͤ�:&���	��Or7+<`\\\˘�䃵|x�C�Ǝ�8��qe��>R�'������1:/v�M�\HY?Fo8Φ�A�A�N
J�C=��=t53��/��Q鎼�EeiS7�B^ގ_�p�c����	H����ɷ��Z��䋦gV�諣?yv�	p��M�$U弬����q9�ɣ�\
�+G�I֛_۲l�e=o���g���5__��2D3Ċɂ$��a�0&�z1M��o���">�P��ז.�l�Sȹ�<#*����4t�������z]��VޟA{�#C�����C����t+#x�� Q�Pe@���CζJ0�u��h?)_)-�S�����@�L��=y �=����{����˩��������6��[�ѻ@fx�Z2�3�&$OȪ���R�Ծ��6i1 Q!���7��U��P���b�ҲF�&x�	��k���9��C����޶��3<#v�=�>�&��5�K	kUl�3��˪�霙0o1�i�C=�e:\����"���u=� �5E���s� ���Q�C�|���w(eiA���,���\���bF[!A����Sfģ�L�-}�
g����`��m���􉢫�m5Yf�e��\|B��i(��Τ����^�;l�Yl2L˥w���
�]�.���lۭԳ6�gjD��.�"��S�s�,���3��o��*�u	���� ��wm�����@�`WI����0N�O��j^�H�����P�7�Ŕ�:6���"�H��ʹ�z��(�.US1�%�h�d9��c�#�H�Ia���)����w�75��,�����5��R	A��w���c�����PbV!�Xi����;pj��A����K!e��ֱ���M����~�in>4���`4���+Yj!;��HE�vgT�x�\p�f��_���O� EbT����А�y�̬V��1�j�yE���QƑ+�}f��J#%s(3;=�x>�	�!V�������tt �){T�@�[���"ͤ��Ca��<"L}nb�8��+E���rI���*	�x�n`$�5ʷ��\^2Ԣ����Y�/J^>9I�_�L��tt�����s�������o]������+������X!�0��& e�"�x^�C=�I�l����$i��/0�C���z����w4)��]J}G��=���wb�$�������'L�{�Čg+�S'��څ�����w<؜�K+��0��`�d!"���J����ٌ��w�v���_+lԆ�"����ѓ���YyZI`�'Lnǲ� I��i3�U>�)O4�gx��;q�����L7:�ī�E໱�Sq���ݥ�sN�穚�E��E��w��Eg��|�'��q�'`R=M05���������!�7|�*�%`%�pwa��ÌH[�PT���x��&�'�w6�x�3�eq�yxNZ��Dt�L�k@��L��d��m����z����u�c�sŁT��a�hM�3$��)�@��\u����B��b��a��Y~0�F+2�D�]Dy���S��/
]V1냔V�pY��?:߱�k���W�o���Þ�d��`�y|^*e��s~����2�k��B�bm]�=&zăA�kueM����0�$ʒ�j��SnX�/����b����㑔�`�uχ���L�^����IE�02��F�v|�C�T��5lu�ɒq�f�e�(\�Bu�/=��1��G
��t@�=�Ģ�6&�Q�<�Yj������m��8�m_|��;��q�/C�db�'��֑�#+��Fe/�B�5.B
|�i�i�