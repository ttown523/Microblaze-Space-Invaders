XlxV64EB    5185    1230I��P=`�O緼����ʙ�T����7ڻ��^�p�*���h1-�rc�s�
���%w[�>m�;�.��Bl��%�ii�q��nKo��@gJ_�ƪK��w
��A��� �{��<* Ko��򇄣H6��@裌~�@������M�v�����f�ß,�L���Ի<߹��� ����6k�¡���6�S��W|B�Ot���qo.�Lհg�����痖�-��U��!V����J�����q����b�-���Q��#'߼��Y{O=K .��~|
��$o��5�fq����9���є�<"���l� �Z{1��, ��]�e�jꟐ�j�D�׹m��5oS�gf�R��"|�%$5��0�&��?C;�6���c#M��E�Ĝ�1:	�X�����U�@�A?>�e��͑C[���̉O�n4��l857�>��F�>_;���8���N�OT�?8F�Y�j�L�K��~2|�y���-��l���I�|ɐ�� �*�Օ���>$U���5�=4nb�v�
5�$��5����nٛ�B[���M
��� .�~�C��!�3x��;j�r�.�e�Q�9�Oѷ~�M�gO��T�:ڶz�+J�s9h޷��8��!�n'�}~�xĂ�W�-2:+j�v�|G$��I��P����?��
�&*�Gn+��g�q�HT��|�%�i���������rV���R}rzK���D҆{��(��B�A�宜5�T^��N��C�L)ij�R[+d5F��e^���@���ҙ�G>�l=�E�_����%p��jy�續��&�پ_��ttر���Ń�6��j�'�	@#�ոǎR�Y�PQ�@��]OYט-��-�-,�	5!�h'iur�!����������[N��I�?�@Y�u2?_ ��jE�b�>�>��>-�q8~�Q��w�[a��3i�4_�n����cF���˕d���Kɨ�vzU����E(IUE��[��-݇��/Q�&(�y��C��ӵ���X�v��Z�E��׳1���yW��������)��A�F�>O�{z�5�'��t��Ί~M��q�e��e�E:�vRQ�9������[w�%�ƥ�P2��_�yԷ�IG��X�f���Cf1�%���&��t��~4,��^�S��L:x���h�s�.=��14����m{�3��g�`�Z}��*�bcP��:,5��_ot�~K����J���J�O���Al��~'PC~���%� �
	t��5Ɏ]զ6N���ٽ;���9��R��r����_�O����N|m�bR,�� $�$4�1iP��uy���$�~��_���A9��x)�j�D��l�ݖ��Bw`-vxE�WX���u���A����n֢hY�rv�!� #Iso^�m�c�6�<퇓�BZ  �79ƪ�'J�=���F�t�ʰ��ߓ�O�`/ў����Ո��:틵��Ų,��/5��O�XB�#�-P��_[8^(��ףuI��~��<@�I�_o�@�i�Ǹ��cE�ǿ��a�r�2���>�2�G\įss6̎�����)�n�[#
�,�}J؋�&/oH�ْl`G\��ڷ�o^]N���3eyT�?� ��ci�
�
��V���?5�T�h(T\H��	��wq��п~li�oЁR���ىm�{�W\"sI�Ƹ����)%9';�^�ȝ*B$fj@	���
\6P� �pjZ��~�ۋ�v��	��ᇅ����2��+���-��Y�ׂK W�f;Ȣ�:eR�S	a�Qy�b���m��tʉ�y@�����D
��db�tX_$��]U'�F�7����CHk(�8ʆS��]T�� ���?�ۻQ஠'����x�B��EQI1�������;�GXҥ�ޟdWrk'�s,:�����`��T"pM
Do��bI_k�sA@2}U�k���V��3�g�J:�}�#	���e~��'�Ș�BӐ���K�a���2�T71�����j��������� �ǌJ��#�@��xѧ�.�7�)��'�]"�wY�A��+�3�(�/[���@����hy�k�I�]�=7�瓙�bcqKqA�$�!%ư�HV ����d��f�5����D5(�"�$"=)�dGwQ6�$���=6E.CAۙ�B�����/���#nB�d:�:p��4�J_ ��_9��N���o��Tܝ�N?�1]/���Ohݣ�#55�_F���SJ��m?����:�L�� Tv�D�o�����ŷ�>µ�^��j/>1��"���Fv���sO�?��0��c�����qt���X�FW�B)ś��ߨ�%fn�~��}#�k�L��3zȫ��Q��B�7�>���K�����%���D1_`����oXٛψR�*Q�1Q�h���E��-H%���rE�4����g�l� 4�/&g�	yk�R�>T�'�����<`Hy�fC��4g0P3�R�߼���ͥ�>�����"��"K7yd �2�I��g��i���T��̚�`�l����P&ݬ�s��ɉ�X+wH�����]p�&s����6�i���@��-������]��UQ����c��t����V|Hv����4܇$9�a�dZ �ڷ��:����߀�[��F���[	8� ,O�s�	_��hV/�r�?���qL�������W��r�����Ζ��ڔrL�����y8���_=�.��B�5[&G���©w�:�Y}��,��� ,"a':�búd*��/=�ǻ�B��m��,�N���]^R��9������t3T��=����)D,X�
��5��W�L����h.��_�^*.kO� -I�E+N0H?�Sj�}�r�Ôa�q4�h��%�W�֞�f�b�Q���2������u`\h�V�)��h�gP,~�g2j	�O���݋tj-C��X����~��!�������.+%#��:̶�$k��f�l�$�ꥼ�ܳH��aF��ՠ�k�*L�pX]�q�Q/�a:�-D��Q&�&�9#�5��M��JuI�5�� ��8P5�%S%�i���k��oQ�%S/%����<h\��ҭy�\���a��@v��^������:@g0l�t0X|��x�zf �����H�v�D%f�?�{�/�8X���0ngü��>x�k_�yrN�K-����x,��<\��q�8�O����}26y2�y�A���*}H�K��xt�&�	�5H��,}��
.�(��?_*�t�)888�u�b��
]/�U2rh���|~C4N<o����`�澀�Z��W-�+�H\uzǵe#H�R��m�$'�D�T�r��e+Û�NJ�aX�u�
�3�[�0�ٷ�3���b�2~z,��u3�WR�S+K1}
7ߠkM����Q�*Wu,I(at����U wE�<��Ƃ���(7�T9#6j�'��Kc��u�[���@s��hm�ע|/c�	�a�^�Q.1L�6�t�ڦBT��k7�:��9��A���&��	=��V��l�p�?i�b8�=,�Amr��BP7iѳ��zWR`m���S�a<� �{�e�h�=������Y$�5!���k�A&Am��\�T�
�����S\g����1��is`��<�ky���PLڪ�e���|u�d����M7eBM�T���;�G�3��Rm�:�=�T���,������i<��6!p/L����8��)�׎Qbqb�]�H������(�X4e����*��'s��e�5�^3�kjc"�T���1����8��N�m'����P�P?���c>|+����M�ކ�2-����4��7���%���^lp�'	�v��dG�Xm���+*-Nxx��:s8��3<.�UH�V���<��2�N�ڌ&�� I�W#u�[����\��B-��8st�<�}_ƿ�/�GBlZ���6?��TȎ_/���CJe�:�_�k>"%YW�=w���F�E��B[�X�B�5n�L�a��-^�Lɒ�c+�K�^��r'84�s(��6<��KdC���޹��L�QAp��������0"*w_�;)�m�ҽw�,�֠�C෧�7e�t��펋�*h�_D@Ќ, ��uo���10=Z�#�ʻ�h#l\�.+�q�$Ʋ�[�c6U�͢U�Ҙn<�U�),��co#Q�d��O�Z,�h�t&v�o.��a�9�,��Y:k����p$��� �w��͘��fFh���(s�G8�Z�2I�4BF��c��[P'��+7���_�د8NBag*�.��%�0��e�_�8�>̑䭙5WD�b��H��<�Y��4��N=�s��4�-�i�J��o�~p�Y�CXA��BQ���B�_�_��bR�	�#�<�q����=�P�8�+7KXj$�����%d��L�y�Nzt�io��cF�I6����q	om���3���E>����%_ƽ�B��+�c���`��
���gָ���G���7�CB��ڼS۫#61����1o�w���;h�g{en�vo�,�6g-.�bx�dDbE=�ᖍ�r<������
