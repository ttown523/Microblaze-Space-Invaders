XlxV64EB    3ff9    1100�g
@0�!g�@�1@�QiݤTǋV���@38_V�s�Atn:e�<w��:�uU:�N�^����Q��Z^�(�#v-�ďLe>�E�L;-H�l�/o $��k�Y��MsC2��1��TRz�^Z����W�u����:R��͍��0d1�O���-q�Y��
a��������|'���� �>1�����~5o����3��3���2?��e^R�=��	�;�r."@��:�n�5c��6�CQ�W��W�ao�M=]���>�[O���ˀG|�B���qB��$f����G����?�3X55���TGTK  ؈D懭A�KX��G:���S�Rp�.�J�AXO߹��-�~4zͳ�����r���;�zN����M�*�!EJ��kP��m0�a;M��E@$�꜑x�J����:�Y���g�^��Ą{2��k��E-���F�s� �Pk���T^I�?����b��5;�d��w�'~z6<�4��5.�xd�s�.��Z17e��4�I�4�D������2=P�~�Ms��>�HBT�\߾������[lm��Mg���W�\,F(�#�����̓��}���zw�.���������Ъ=�~�����7[9׺���G8K�����!�}��Wv���{n��]\�x�h#�Z%�1i*�%�C˧�h�r>�9���CT��Aͅ����JI�R�7)7�ui���#e��s��� 3
�6��VM8��%-�c�]ϼW��&�/لK�ڱ�X!�dY(3~Ŷ���b��Lg%s8�%�t��U�g�I��dc
t11�跄ߐ����/����0�/�eM���g�����x[�yꞗ¸3����)�C&�M[@�����:�h� 	_��"B�s�pVb7�w8P���]�=%%�I���k�x���o<چ�2���ȟ��GR�Ѱx�[0UkZGO�|����3�!v����5]��Kf��Ǚ�'%|�d�%z��]����h��"��� /��v���FAf����lݛ�|"�~�<,��/�(ZR�ay�ʟ�v��m�+�~���"\&�F�%���d�xY�C/v$��e5��/��,L[�q�8��Eik�a�`�NH��S�ᭈ#�/�"�U�c��Eg��̈���$q4+�B�)����tO���o��D��k%<n�u�g�H�+w�C�������@ɚ�b�b,8=�Aȁ՘�l�]Fd�Ԡ/w�KV)6@/ 3XkVxHW�E���P�m\9/��=�s���/^̸x�,�#�6�R9�s[�+�R�c�ص�f�� ��l��#`"�)�^�?�1'�����tPn�b�~ou����j.AߨW���64���ȍ,��/��i�,ՠң�KB��}����n�'��o��{y$'A�(�ap�A�20�~Ԑ��Ja��m�P�Ia����
�(]�����o�!�����x�3��K� ���+��[mD��N�@-�����̥���n��9p'I��59+r0TM��JFLk˗]�}wA��mN��Ξ�w�`� �%�A�o2(fM���d�(2�"]`:�/S���}���1��JL�@ @���G�p�/�}\p�$"&����Jk�(- bK`�Z����Oj?�@M�S��Z!k΢��N���X��bgm ���������M�{Y�s��?��ST�R�����A��=>a3�\Eԩ�� _\Fn��I�2��M�oS���='�������J�P��uF�k�4fԤe��%"�����-����Sԛ�z��[�;G$�`�6�3
����I�w��+!�AR!���m����,��8	�}J2i�t)�n�6�`ڎ�2_�>�N������j^S�M�+���E!��lY�r�l�-�{��t즄��*N���,���3Rk�7�=S7E�p�R��V-�#���\)�-t˨ɘX����!����9u`n���㈸�����W��@F��咹��W��S|JI�(5�eg�����8���Ol��9���_�T�?�dc�x���C��
sm��w�c�!TTf0���-�\!OW#�� (����l*�<�H!P��Ra.t�8�� �\ p,	�op�����ˡ|��>��ug�Z� Y]��DWTn��g�e����i��{�h�*b��q>i6OGη�X�������t��*5�P�Wo=*�����? ��|�g�{t5_�WR&��,Zz����[
����H��P[a���XA|�Hݵ\k���*���cR��a}��5)�2���t׷�],;=-�^�SrHN<�nQ䊥�(@�-���׎����Uo����j-��������延U�INDM�M�A�ڋ�t����ݸG�W0��2��w.h��		�r�;���z�h#0{�k;@��ٸ��\�+y��x��)�:�K
�l�Q�e�����:Ƞ�
r�f�(�Ϻi�_RoN����K�8�'}�S�C�Y�aJ����M{5�ac�PhݮF�T�ľL���\ ���+`�QɍT�R���)��?����l�ՊB�$���+���~������l�T�f×(�J�At�	�\}+�3A��̌w]�)k"qzj��e������&��) p��yLcR�3�r�J��S_����yo���y]�@�˺�����u��8�#X�Z�P�����{���\��l���y˶�����%�G-i� !w뀸�P�_�I�O�'<�g�"����~ȷ�!��y[ỹ*�����%'4�'V����`$�|��U�(8G}a�b�.N�y��Zɨ�O!�R��L�k���h�Ϲ!Pw� ��$��DA��"i�&Wbm���ꎐ D#jk^�����L����p��b������*N��Cb���Nn� �!��n4��7=�}l�Hgf���$LU���ށf�:���|�A����m�҄�Y��E �_�O'�Mk���	��e�^�t��%'��=��,jPx<SG�����[u�`]Ma�B@W��->d� ���L�(�<�ʃM��%�ζ(X�� h���W��4�@^3 c�2U@�<�9c��N�1NR�k#�`y��ƜȎ|����G�v�dI�q%j4`\�֓&�朱�.���S�#������R���;c�7g޽q;~:�$IX�)�J�՞/!�{y6� �J�R�Y�����������3�x|�3�&�A�r���;M��)���gE��7[�C�-d����I�)zs�e1�g���R�d=�������I,Z��2k���?�l�2H�I��������Gn�pE��?�u���u��?��?8�r���#�:1��ǧ�cojp�,��ַ2
�sS�2���	FGK��,%��D<�j�i��������)�T+e�U?�)�x�l�����)����?'[g�6�>ʭO��O<�٦1G0�Уm�ʙ�qW�o� �+g�K0��bP�<sN�Y<TzҾ�� �� m0א�1�(����N]L�@���2���RLj�hh��p]�K?�(�gd���y&]u.HN!l!�����۟1-:�8�s?V
�T�(�#��|?���\Z�nЉQ&�o��Uջ�'�bJ�̸~;خ���P%��'=8��Y��;���tݶ&��h�}%U�� /gM,���.p�0jw�?"-7u�["��w8Ad#���t��_Qt,VE=�k� ��;4FHW��1b�w�݌/mfm�X�#�]��Fu���wɹ�2YX�^�;���B����Ƿ/rX��q��[�o�#�Y^�O���T�0�=bo]�N&F�62�����p��iYNU�Z�J�@��*VJ�Dx�Egh�#�uk�Z�,�5��:Q,k'�N�]�c�)Ki��W(��	���ۧ��JDE!�p�j&҂S*6c��=�ps��蔮PK�[s��.��f����M�I�R�s��b|Xװ[��d���?�k���=\�iulV��'��z
-��p��	�_kd�������h�l��֢Y@d2��e�,w�)t���f��M:�R}�����̉C���v/��A�>�Re�A)YP�u�%kV�$�HFt������������ _���Kr����:��V���M�I�@7s�^�3a��Bw���Q�%EMt�!.v��;�|��R]�	�+�R���	t^��4ܕ��V�s:e� �z�;��QV.�e�i�m����T�؃sהwsYd#yGN@I/ N�	#�U�N	�a �y_Gѷ0�f�uc
�T�H�f
	�Z�p�l{P�b�6