XlxV64EB    244c     c00C-i+��wѐ$�P�!vU]F�_w>�ԢC�MǼ�<��
�	�E�*�2�p����z%�Kh|t��+�E�&�*wgl`�%���`oA�u��.[3h�#�8�)n>�:�ٓX ��c��9%XL��2
��+�;�������j;�(�VE��y8��Λn�j�U$���ǢS/#�*��u�~AjB:�����h:�~J{b<ٮ:�f]n�1�i*��s+M����م�6�O�����>+��;����!�qݏ���$����yi!]xl�3�6�3O���v�m=�3z��]���L��>�K��B� ���H���%�)�F�8�B���y��87����������k�n��H=ܒk^�0B���\l�,���KV9��_��,\w�m�f�%Ѝ��!o���c�@���]2���;�:�74/;h}M��Q}�����Aʘ���e.wķ���>�z��L-���� ��"��x�*����+����r�����Xf���']X:�K�-,��9b;�{����\�i#�!��-�'�	���@	T=��
�/К1�uX������K#G�g�CE�;�@���P -���e���k�FF�lK��F�7��.�h�����y�]>��#�}�R�i�������A���	�����e��8��1��K�,x�w�A�n��ظ���ҝ���^j��2@?���B|W��A$�� W���r�%���F��x��AC�]�6��GP���(w�H&�P!�s��6r?����j��m���,@��@R�(� ����Gb����@�a!B%֓]���4 �԰`�����9z�,>bm��';�Z� ��{F�K��'p���(}Q6����M3:��#��>80���5��?��/�52�������]L\�����b���|����dQ�,��c�Ker��L�$N�h���UM��vYo���z(�,D_T�� 1��k�>�Ԏ�8$&�UN�%`.�[6�,GN������E����l������Y�w!w`qSB� ����Ȣ�4�N��ۀ������5֩S7���Lܣ5��*����LX�&;d�Sb� �-��ҋ�l@\m�n,-�ϴ����az���=�t�AvQA���]��gM".��zON��H�×	fN�ZZ�f�2�n��Qf��lllh�mn�HgYx��v�A$*�Oέ���<8��0��`�졃leun���X_���������`sL���e�W"��a(kV+�B*�R��)Ć�M����N#�(:7�ma5vG��������B����x���(*|ъ�k�c�h��Cs3h#'b�#F���て����
}��en�f�E<Z��+��a��ѱZS	�6�[��UaF�Br�rB���fԏ=�B�-S"pO~07�����F��JC{ݼG����bޓ�w3�c7�gLL���%{�Ώ>\'�w��Tc�A��-�t�+R)��\x�KE��3Zn�k7�������wr�*��K��+.Gz��𡢝&Cw�/���0� `�#-/NP��v��P-� ��폛Q���[Ϗc��_��g�C����L{�-*U?�B������� ��)�:�$Ob-*��z��@/���3�a��L�cج5 9-.� Bq�@�џ9�~��6�d�MSL�r%�62��>4�F�J�p1Q����&����7Ӳ�=�P��j��dL�>OG�9i~�P<�E�LB�HO욧�O��������Hhi.ޮ����<��}B�q��t�uLȱ����9���9[7�~�n���3��$���?y�^�$�J"��`�'�
���i-�$����Pd��~����e����Y���?��U+�)]�f�EK�%v��c4� Xm���-Q=�zhs�&�Q�J����A|}�tP�bd��Fjz���A$6t7���������T\�+<�7�DD��5��>�g������'���r�D�,Oh��D����2�ܞ��[��3��n�%U �����&!@���Jd_�8��V,��P64qbu��y���2 Cj�_zC<�]}��a��&��TDo�����?d���+���)@��dTKU�y��놾 9��s@��f�?�4�ˏ��O���U	n]V-�>�Z���ߩ���	���5+�� ��׬)D�vj{�)�_k���_�Nw�0?��׷�����u�c�X��yY��V���󰡋����^�����s̊�d_��R�DI.�U�Q�w�:�zz��ovv��D��E|�%U��?Ɂ@��É>Y	r�Є:�ֹ���E%Or� �� 	bSJ]u7��zr��B���	0�gV��49>eBs�%@���O���N�N�J����8|���������jT��V"_���0�Q��bqx|5�17��+��@���W�����]i��d�@m{z�����.�<���_�g���Y��=��4%�Q��+�0c��YY�Ze����)�����(�.�DO���M�(|����cwIZG�r@��6;�Rw?����h85��t �f8-�*��*�;�Y��a��5g�l�TȬ�R"�L��xlwn�KCi�\h	��ҫ��>l*�y�ny���81w�[���V����SqF�;16Ȱ�<_(kS�E�l'N���I����%�<�����ļ�"2����Sř�����H���J��.�Ƌ�p�C����h�=@P�#�{��P�P���Ud�׾�����$�/�O�9�~�(���j.��/V���������5��Xn]������r��(��pt�O�ٚJ�f�vD��v��/���r��b�'/ �����%�l�e/� eX�G()��FӇPOxQg~� `UOm���Y3F�+����_���KC�k�J#�]�%@����*~z1�:���j�3�3�h�����������	�p ��;&�lB��֕��w��?s��(��1��M`e �8Ä#��vHU���aȱZn�;"=��