XlxV64EB    32c8     d40@�e�m��=4%�ߵ۹H߸�(��O�� m7,2�\�n5��s���&��ZJ5KH�d[h�5����72��@�9Py�З�84�M�nH��M��Y((;�7��h6����:	���3��J�N@U�����|��]V|''��;��֛�!��n�h)�o��B7 �����d}Г7�.���켶`��ٴ{��U�pGM�<��:+d�`Q�k�־þ�Rf~���8���O�B]����W�eONa��5̯�=k���h�b����Q2b:��Ô�͆�>�n��kK�)<3�ŒJ���],���0z�m��� �X\�ܔ��a�^o��K|�"������-�T�����79�?����� �ԗS�@p������o�j�������h���}�>y
���ݨ!���f�ե�U�䃥4}��߈p�u��◽o��:Ğ	���ZǛ8�+MVR�h.s-!N�k�K˒/�\\��]�Zb)���.�b��Z�����H�����(��Y��$J��o�s"�l��:�:0���Ow��J?����Z	`�bH�lN���"�bjHDT�F�-.�����b�9n6�VXn��Y���`V)�����_B��N#3�5�Q�_~��h��*3?y�u�^��!-���&v�YX�*�S��<s���@NXr�
7_�/������|Pbcδ�0a">ڊ{�H�SY��-�#��+̌�ؾ"���^��͌�\s/�v����ZTg0���o��S��4H:���uSǴ�H	}Z�څ�Wr<l���1���g�k��b�0�W:�v)�'��DR��H�~3;�x���]�2A�k��:2LV옟���; u-Ĝ��IlZ��W�d��|8��4+h���e�J�_�����ā�1p�&��rY���f��s���.������h�Va$M�v$߾
x������>[b!7l#2v8���m/��Ҕ[��WIw�.&�n���&�I�4�u���I�����R��ԞU��S�=�ٮ�U�u����<���������i���l�Ʌ!�yr�:\����;b*�&�,>A��~H}ӂ���6��Q�}."]��([�M����� �/8d���7��A%&H��)Z����'<2��yiz/wb�\Ȭ�͔��*��K*�X�y�-����|	�N:M�I_�;�9~E(R��u���0���i�l�Ğ��0����=-�ḩ���+�n��h�U�p{"6�C�l������{�#�g���[ӥUn�p�	�e�
���R5^`ގ�:P~�YB�d$�yk��D�?�|_�e?���0F�׷�V�U��ʇ�̥۟#2a:X�!�����4�ȍ��A��$�?�DR�}$�(�m��r��Y��ٰ�6FCg5J�%�3.+@e_�k���|��e��/���+�l��2T���\�f�+�� ��������BH����L�"��b!A�h����a(emUk��������}H|�Y�_;�.�ƭ��ߡ��(��w��'H��*�n;��S0�@��{�i�6D��rMl2Θ��o*���hY��H���,T�����p�)�b���h�ΐ���pP�Yh��w���~�C��bN�9J�������I[�;K^�[g{N⼚�?)��J����>�b�������w������|�����a��=kɁev�Y�rm�@
�چ��k��@`��W&Na�n��=�h\ <�US�����o���SY}[Sʆ�yu��"UДj�1[��^;�t#�T�F1hXa�c���<7�
p��L=�k�ֽ!�� �-����_덆��_\AY�Z�NϚ˴�D�臧���Z6�QD�|�Y�#�\�AO��[��{�s1�&N����M�5	t��ά� �dg��u-�d�5���~����^����`��c�;/"v��`ܲMxf�;�_x�;��M��ԓ���Z?�Z2�A,h4�lIw�d�Y�}m�z&�џ{/V��M���LJ
F��:�����Т3`���&(�c�ö@.+g�) Ɣ����W���m����i�.�<�����J�<N�Tva�7I�iN�s���x^g��_���F��1n�v���O�<߃!PK�љ��o),O���LǱ��ڶ"xD����b�o��O}6�����z���̋��irT���q2�c�ghk~��J;�}t����*�GE�/���L=7.�RM���!&�j�b�x�/�E�E�q��g]fc�1��D�BE\L���J�A���i���N��v_���n��������f�S23�X�^;�F�Q�.5S#3p���H���'/���P�kӵg*">��ԀF�%Ty c8�EXK�d��.z���|��]_J��9Y��sq�g��σ@�kܩ�|T�̗�ŤU�Z��y3O��f�_]u3O��S(<�K�������g�� �D(���V�e�s	��w���W�2w�Ml�����ԞM�=����K�ק�����l�C�s$OY'!nD��弶c������z����Z,���Ǒ�)d�3�\��Xcg�����o?�4��aQ#]�J����LJ��0�{�׃���dmaH�*v+��dx]$�f�i�|;]r�A��dywټ�����~�q��ُ"^*kR��~ i��D~���8��(���>�;Vɾ�hi�4��9���6ځ1H����f���"C�R��M����y�
����i� .X�ϲ��)F�@�H��'�>>j��������LB��Y׺�㣓n��aD���/� ��\ )"+��扬!��Æ8ނD]�T��9����&f�\;X	�UW�f��fӑ���g�S ]��@X���i���]�2�ٿ�&cR�`�����5���6�i7����-�����d���I��vL���Φyn�+:x�2��X�(�ά��t<,m~����Q$1��Xid���@�2�8~>o�+GV�3<�ȝ�����ZI������6�ȹ���ۊ�5�ǿ3�6/t��b�]W��T4�^��̠S��PzΒRя��J�� �H�и��ȥ��Rk�Z��ܕW>d��E�v3��'Q'���ӈ�.�4h����{����q�f��a�Xy��ڈ��sa	w��O�T�<s�qK�f��,���ׅH%ǥ� �I��ǿm�gk���.���IYm��x*)�������@��-:��^sO����6�-]�\N&�g�n��ho�{|*�fE��h@h�f1�/ܮL�l�{�mu;j�&9G�D^0�6U~-�'��j��/�l�h|[����C���z�=e*