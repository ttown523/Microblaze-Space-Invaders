XlxV64EB    25be     bc0�&H���1Σ��52���O�1��a��(�X�)��Z���e�+�ܶD���﫸�Z3�;ϡp��;s�h�1{1I�+am:����AA�_���N�P�a#;g���z+�M�ur�]�� �K�n�E�r*�=�M�O[��7�]f���[�Q-�o�T�J)z5	��7�h����u�§3��S���0P������e���V�9�&�D6F4�Z]"��(�N��Z^�{�In����p�3]Z��l��
*��+]VU�H��	ق�>��,���!iR(��fP�G�']{vᢀ�	��V���K�3�	G�l"��\�v����0��Y��f��'��
|��N�n�	��T�G��H�f��9�v��8a��z��w[�����2}GEj����5nw�#;yL�ͫ���'j��x��G_�%+�\��o�,�f̧{T'�+���dW���/�9�~z��f���z�\���I�(�-�k�q�GI�y�����!�s�so�%"ѓlS���,������ 6���Xc�"�A,�D�P�ٿ �7�@�rW�^D�~��H�r\ �~�Z���>B��(���ʹF|��y;̌Ȥ��~�U�po�q��v1Q�8/��ī.�O���Y��V6ޘ�/�u�s�����7��" ��Pu�[�>h������l��v����lK�$]`�U����v"~����ml���!�B=���4�nP��|-j~X����J �g���W�)��zu�쾩6�m0�*�_�${�:Rt�-�*��ҹSCa�ǲ�uvx��"������RJ}��
���4���NX&�.�f/��=��xma�_�Xwf)e�8�X��܂��z䧝�P�~���0���zS�H�6�Gd��E��L@;��׉��<�b��[�b�
.X���hx�5$dզ�7L�ѻtD0Vw�q�p{ן�G$�[C�����.��|2�u������	#]D���GG��/�U�M�A��(;��+cd�Sϯlɒ����͙�0h�-���d)�~��4�{wN']���2&���%e����eє���+�������})�{��4�",^�9�04�\�Қ�oo?��<귮IU�!��W�Z��gV�پ�^���W�$�L�E�Ƭ��g!hnw96��ܸoD)�
/��ͨ���I�Kf��J˕<q�A4fT64��~����'���v5E�ݑN ���v<0 |�l���e�сm�I������g&��P�p��8�*���A���i��󎓾'F�ߒ^b7:�xY��v��-k<ȇCU��F�@���!�r4��x�W�>���[#�f/�TQu��:��Eh���U{�>�s�=���!;U�`�"�ж=���\$
\��J�ſѺs��ȫ�}�ӑ���0����G{���HJH��5'��]�v��Խ����9p
 �m�S��	?��RM�y!�u^���Ļ�'\�rL�1=/����'2A�Fw��R��}t�J~��ܿ�O9c���}V���S�E���󨽺d�����&���S�}��HI31L�Xե�C7��k��pH)%����>tB�׃�g.�æ���Ψ��{���g�zC:Wi��y2ItI�e,�k��?��c}31L�:��2E�.0�+���K�C�g��{�:x_��r&� {jɍ%��qc�q�{��s8��`{���xd�S�������P4"ÚA!��q���2W`ym�G���Nq�t�cŵ�T���/�Q\�--)�ڨ���Fd�~�P��[:Z�\���P�ג��]��VFsI��G��Ĉ>�қ�����`�Z�N�\��ޡ/,2p���|>i��A��}��9" ���7I�s���TlwYK]C�
����&�����B����n�m����뿲�;"�ڡًz��H)��9�1�rs�I��_[�eԝ�&�u%��8��ҙ��p=�|�,�F���W��L��;)1 �9�����䄃I���ﮃx�Iޖ$#z��xו��^�x?j�-��i��Q��I�E��DN4�?��Y��;Y�|���l�
�y��;������x���9��)D�ߢ��Z�~c'F�V��ӻ�ʦ%��(�F5J�	�~�F{��I�>R뤆�������?@2����}��V%�#��-�$�iK�TpOa����܅7v&>̭s
�Ts}�	A[Μ�Go���\]R%�I��U��b�=��vY�����������;bQ��l���ǘ'S����x�yi�����Ҩ�s��#������;���H�Ǭ�̫�ܪ�������G��QJa�o݀�G�ol������[҆/�=��B5R-����5�}�~Jo
�U���J���o�=]��hSX:�8��sH�e��u;R^n�="����xRԮ��B�;��_�Em�
�� UaO�?�Χ���[��B�-��,�����\��R=�͂VQ�S��W�My�&��{ipg��{���:D,Aˁ'������5Gvq6�s�Kr�D��Z/���ލ�nD�xs���X"�9����5��|K@2D��Gf�=�l��f˒YD'��D�	��Z�s��YA۾`�9'��F���Y�׻��g��mk{W���֠�G��`�����'��~,%_W�!�-1 r4��(��K�\Z h������؋����Y�q���D>װB��5�s��I_��g�Jٲ��jեL�7Rܓ���f����'_���etX6�M�\��>6��mtx��IbbQ�4]������6� ��f.�}p�Ֆ��h�X(�T�4K�{e�vd[�(�h
!�V�@�w��� �s� }\Y�v{����@�����2����Ia�]�d� x�d &�?�ʥ��V�������=����7���7�
\�N����W�&=���z�X�xƲg�a�D?��٧v��hA�i9Ez��8
