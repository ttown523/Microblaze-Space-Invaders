XlxV64EB    7a24    1a20R�)�<��55ɯ�aJ��_������C��R��.a�?c��`����o0	��
�A���؜��ຕ���F$�˟>�� N��dP=�9OH��B)c���`a,�%����z��	\d	��~Z�C�*}���S�O��\to�lZG�`i8=�cG�"%��c�?m�	����y8o�!��H>�*�/����xiy�G�Ǜ7!	�PD�>캰(�����I�;v�7�!�k����4��5������~����R7��(��~���t�s x$Z�@�[=�+J}�F�����*Z��~���!��WU9�$�Kj�=����ٚ!ht������8Т��F���Ęx�iR����|Q�Խ���|�Ņ�QMCR�_�?�oi$��; L�^�[��^����>���������\V��qXc���,�� 	�@� ՚L,Ѐo�M���=�$1e)$m *�"��~�ܚ�M��z��/8�I���d��p�`�z�U��C���3����v����ml�.MP�֕��2��\_��gّ�K�v�^���D����o3�>���@�����6ԥ?�`g��j�n*1i��:_vP�����pW���,b�QI�j�vM]�+��e�*��S/x�pP�S$�I!û�0f� ckRFd�^ȇi��@UW����;�"�O���?��Ü:_��ɇ������#���W�h���E�F�V��M��S��O��0�t�qǸ&��7֦���泒��n�	���u���G��y�� p�P�/��Z����E�� D؃!�"޻��X���f����X��%�F���԰�O\�� ��5x�J/�Od���ttwl��9̺s�&�VT�G���ۃ�['�m*�ѱ��a���u�,�����ǃ���Q�L_Y=�Z�i{^ԝ��C��zќQׁٲr(S��Y�:�ֽ�U��h!c�HmY����xŴ�꙱��1ߗ�Y�;�<�cB��@:�����6I����%[�O<T߬�C+�t
���,#:�4��D�%���0��@�=��<�\si��[oif����O�N�-�C��ab/<u%'�N�����ap�`��b�[u���@sD��J���f2�j�7��2��#���?/r�12�Z���l�M�J����>� c���3b�'�꿤٘���@�}sG��ߧ*�΃|��Eat�"ӏ�t8*��[IRݏh��4ܛ�H�@��/!������g��iU}�d�گ���->T���|PW���§����>m�z1���Z�u\>CT�<��"D��+*�^�t��v�d,k��t��<|���W\�s��L�5�m��21���z8?\����vXQ���T�xx��F�-\�i� ���:�B�$s���d�i#�M��"��\��\c��^�)��M�
&izԡxt�s�&�1���Ec3�`$���3ȭT��ȪIxR�H�Eh�[i���@d;(%3��w(�C�L#�+e&�Ї9P�0>�����Z,����˭�t{g����zI��z��f\%3�i0:��y@Y3vk�&�G5�e�^8����[���K]��B����;oHyPr(���JN-r�T���ʼd&�cջ�iX�|�8�9�~��SA�ڸ~��.�3W�]�ѓڳ��K1���M��7'��e��;��<�ߊ�'"�L}7�}�C���t�G߳����߾5v�0!��������asn���#yW�
���t7�~n=��Ǒ*���I�ڏT"����#4[ïut x���c�]=�9�u�w���p��� �QI��D�gQ f�b!�F�ǐ�Rroz����'⻒�j��H��wD
ټ�<ߏ� K,�-<�#�F�"��6��"�RZ����>��wkSEn@�0��:�#1������W,W�%�v}�<![
���?)'2��[�������;)��s��������V��"�qc�`0��\�9�r\{a��m��7+�uv�֚�rg����A�������rH�D�$?REJ	��|<��ka²�@��D&^���f�+�}�4�`ڸ�QڃލUp ���b�Nf��-��p�eM񄬣�o�_��x�ޱ����l�mv{V�z�\���vc���U��J���hA�ު�Dk�G��	���:m���23@�P�����yY��(o� ~��e�O���A������On5��bY�J��b��TG���P����v�f����s}�.3k<����"�0-J�r�"+n� ��<�����Z��K����4n�d+�8{���J� 8������@5gKJN1����m�cB!Y��=#G�LxS#k��IO�~��Z2�Zc���Ez'����0j�>[�u�ý�iX�ܟ|7(>����܇�����9��.���>-��5���(x&�M�(i�b�~3w��ſ݀�Ug�n��äT8�Q��U�"�i�G�!��̾_�6��^��˰�d�<1�Yzz��z8j~(X�$������w��}�
5$;Y�	0�r� ���)�rvB%��F�2/?�G�׻�N�*�)�$��<W�Y0+���W_�t�*Wk�.�b��f
{��P���c���&�Ci]��É�<:�Q 9�kR[�8�1��Q�e�tR)v�kS�X?�V<�'���+y�7�p�$R5�O�n��{F@V�n�U	���?�"*S�����01�0)�E �`e���5����@�c���&
�^UU���^Z�l���>B������ŗS�j.�O�F�l�;����lQ��⏱����꺇����F�%Ty�K�������+���, 6!�[~�#�E�~��frØ��g�w6#0r.�Ԗ~v4e���F�51ݗ���b��Fv1���czt�W�`|0�G� �Ӟ�����:u��A�͊pˍ�>�=��8V���e{w磹F:`c�0<FWda�mJ{�s��c(8Ɛ{B.��s�b�M�V������$��1�%Пp~�[7���y�|�����Ɨ�ew�(}�HY=�E%���_�y�W�h!�@hQ: ��V�e�t*�X�0J�2�>�(�;����v�����*����Κ�r\����?�a	ێg���8�ovr<4��=�F�ߔɥ�Q�u�N��G��Dr��-#�^:Z�C�nm��f��=+���Bxr���!����*��Ӳ��:i:l��m�;BM��nJ3�$$v�j1��˸�Դ��]@�V�E
�3w��!K~�P�Կg+�d��u�T��~JȻ�㜨�Y���ɚ^�>����8�b�ܣ]���;���-;��^q-�x�����$��p'k�)Jȝ)�J+5@c��K[�V���8C��(m'4Z�
�ll!�&z��B^�Y�N
��O��"�R��Z��?ڜMg��i#k-�$	4cP�AX�v3��M}S�*Α���?�cw��m(f��w*^"�<!o�� R�Ҡ7��φ���Ǣ�a�A莏}/val���lC	��?��D���W��Ib��%��^�avc�G���anx7h��	�K���$�?�KY�{\��4��7k�*������e�٧�R\]��d
�/�~w����ªqV��#��mbY^�:+ku�5`}^%y̱�pNW!�~n_W�k'�~���ص�^�s�$��EA��w�@;�Gp��<p���A��>)%��"�˸v�+�ѽk3oD:��y1kd����������Yav:��6dm����v׋���n�k}���>ic�#O�T�U�%Z�ءl���V�PK�_��Y\�oV���������A[�D�^��Mo����	��zڈ0�29��b��5���kphd&Rmv��n�n����s��ʳe$٦pQ?+#���z��zXN�c�N��8��2��I�X��b\���]���LLtZ���)���D� <w��f�<����Dvac�#�c�� �!�RK#a��tZ�-���=��������O�yA&�{���)W�A���/��Ԏо�[��g�rו���sf+;�����<8~qj�w<�M�+���'��7g��6��璡�Y}U����P�3��U����F��f$R�E����i���g�4��k���)T��cF��2�����(�j�αvɓr��B�c���l3��*�����?�[���d9�Ƈ��!�� ��`���X�8++��&����/����Th`d [��4��e5 )]���!�*�)��^e�����笚��d��f7�\�����Z�y3�ڴtE�ۺ x�x���t>��C��z��ASb��4v�%w�^ɕï�Y'_�Arx�妣7h�,j[F�w��S�Ǆ���=-�y�e��"Ĉ���}`��6?P�+���No`��6�����G��
FU����b฽K�̮�:Ω>�'�\�X�$𲑖�`�����"��Vm#zΊA���/ ����7,��#iF�i�)�.?�ȡ"�
�n�u%�VU| �q%I��e������=�.�V4�v��Ǭ��#.�� "�A���.h���+�����A'����Hb�X��3z����B�Uk6�� "��E~lNN#�tIi Ԅ��K�V�'�bʏ8/�o�(��9P���9�3t�]z -�%�Le�`��|��4�I����߱3�ek�_���T�Ȅ�*�Q�� � ��w���V�Am'#�}��n.�cJ��3�8�%����<B��L�����J,r�Ŭ_�U#�d���nx-�����?cw�%u�W�΍�srܿw6��8Tڢ&^1n��6�����(�7���8'��Ə~�n;���� -��:�i0<#��0JZI�Y[Xvr�l��L���D17���s�w����3�g���5O˨�|���q�Q�}��L�8W"{}n���|�����bZ����_��1c��q7K�l�� 웹�?�iZ/W%��ŏ}�uN��$T��vk��5��+���:>��Ng˫�W,/Gy]\��5��`&Z>� ��\�_^BK~�H���x{NID~4C8y[�^#{��J�DY#��h	0�1�'Z>^��9��;3s0_�Z��?Pj�&�M�#�V���ⴗ>gZ4/�F�I#mB��_N/���D��J�w�'=K����!�Z\R㣟����r����j��#��U��=���Ȁ�?*�$0�Ly%ު�l�����,G���>'Y[�)$oT��O����9U���&Հ3�&2ekj�=}�o��~�N�.�w�[�zH0�C����./%]�:'�#˅o 3��}�/<�ٷ�<��[�@Z\lL��?N�G�(�����M���ZO��R����#���u�(���A�	r��2�O%�_~,��/�h ��@����5�vB����`].�:xOש�t���*��� +p�*E� ynMO�"�B��P�I��3�[���8�����C��K�n1��,�t���E4���N�'�"ƆV:9'/�ϕ�н�os!�{.��>�<@טæ5ps>�f�A��r�uD[�����ޫMcr��=]I�$,�eb�!�g��W7Z����1蕹S��C~�kY� ����>��Jfxg��>=���j�LJ�/0�[���X.bnI4)��t"�:��䝼�/�h4UGMXi�G��Y���%	ݠ��,���\^�/xtW�͊3�{��!95#N�PC��x^������K}��r�â��D3!Nf#�b�>���+)$�0z�_�%��C�/c�b�Js�V���T)զ)Frl*��3�Vje��3�����:& ��e��d��¨�5ݝ/�[��oԛ�u�ˤAW�P7��@�pڽ��'	�sQ�I�+"I��$����bL��mo��:�uxd��Z{[�}X��.��VO��H�����?#���U	V�#�S������}��Z�[�l�����〦:X|��~����{��"X��4,C�n|鬭ܪ�srqj�fDڒ"׎eR�j��($]�q�yp\�]�ܸ���I�3�(5��JL2,��z�w�4�������a��3��uW�<�M:Ï�K�G��������N?�ɋב��XX�H��еc����{��*�x���Ȭ���t���!���8����ǘ0�3��ؽFWC�����v9ҏU6�X���P�F,������y����|S�! ;���L��+J�Gƫ�Nd����(2���t!�+;X�'�*�}׃�[��m�ߣ�;CV��o�ȓ�t�Y�x�qJa�;���DC_Z��z1Uĸ�*G;�_��?�Ç�
���!w���(^i�׼��$����4��cuI�*��╃	���]~-e��R;��خ%�,���!N!���E���K�?ր�6�'��p��=.$Hh��Ԇ��[b��+�U��ʩ-�:��V� �f�T&
�Zr�.N\��w��=p��^��� ���ӭ�7�}����w�g�������� ���T�k����^���b}u�GFi�%��	g�9}\�QH�[Q
l�[��	F��F���/$L���O	Y������P�T}������~��ɢ�.�f�P�������oùBq%�~��6r��X�