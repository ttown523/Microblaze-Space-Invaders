XlxV64EB    2b5f     c40<ĘJ~�3��=�D��$M���I���!'u�#������)�A�F���.�G�~p��m�.��ع�!
�� L=G�a��D�f��I�OJ�7BZ�����8<�E��H'I���:~]60�D�L����S��
���XX�=b��ւm12�il�t��L�)@S��º.,�5a.*��y���u��a�*i,����'��9�� �~�]�H1��T\7x���-��3�т�k�����y����s"�����I����Ѿ��=5Uu��n�q���U��+�&�������v�;c/�D!x��73ʱ��7IEm��ܾ�eN�א�$��2/8Ӂ	��)�~) �D,f�nC��dx��Nh��"�m?S=�cQ�ʻ�-F�Y�YB�@e�uձ�9/"ų�)���]\������2%��J�_"<hy!��<&�~�D�(Z�/�7���:.oC\��G1��٤�i	*�oN�dT�%�`��y��s4_x�'���?ʥ��E�j��Fy�D�p����㉰c4��+�#�*�&EV��2?e�1'<��`U��c���	�P��\[H.��S
n�X����9�9͔P�L�m��~w�$��c�w����@-*�����^���g��]�SH���J��]�L�+,x�'�w��>,�+�=��<���������!��8e?�����6�4�`�H=�m��~��Ő�2p�
��6gX�����X�h߫�J�B풍��b�~�����E���Đ6�\�C��G�!���a�)�������)R2${�[4�V������7U��]��TڕЛ0�,�73�VC�����oT)��P�E#�S�=�=(\��?�_��Dx�,0D4|�)�k�5{��D�r��z2A��&�̈́�K�}o~]�0S�'230�q�̃؞���#v�����O9�ƊBM�	 �K]���0V\�O����$2]���X`qYA��>��Y�$M�1(i�$$��  ��t�:#�I��kړ��-��/���갥�ڨ��'��2-�m�IU��9s�<���Q� E�{a��_�ko"k50�����2dҀ9s
.E���B�Ҟ�����'����;4���;j�H�J���=��bƋ�9d�� L;�N֬at	'q�O���P{BF5�)��wt`^P��2���#C�S	���O��?0Z���Rl��dQ*�N�V�1o���1b��o��ұ�Bq��D�����y9���t�����i�v�����}��E)������uyά�=��<B�����]�ܴ�O3d��E��p�0U�JZ����&	n��t:#p0�'�º�k�6� 6=P��ם}�n�7�����L�Mx]r���Ťu��!���g:����(CSvB݀N�~��
�κ �Vk@��vi2(��\Q`���]k4w����T`�9�R��8bx�4���:D!.:��;O�z�)L�Q�]`��d��"gcb(rW\�
혏g����z�ޛ�K����U����LC�ԉ�ex״� zy���Z2j�9�8�.Rw��ˮ�Ag��<�Dm5P4��2ڍ��T��V4���pkE$r}�#F�/ӕ�#E�1Fr �:��J��G:<�7�W�֍������Z�['�ށ����[�CVlh��m9WTVH�V�K?H�|�Ѹۃ�e�i20I{]��I���Œ�����]�݂'�nt8l�����B�r6�	��=2��'���Y"��h�J:E���)X�޶�=��cѯ�5��2<"쑙�K���kh6��a/�U��lCDM<���]D��zM 5�}/
��ɘmIby�^$�,�,��c_ۗe�����,���� ��OS�����Ir�V�OEh!'t���1�8ܠ��nA�Y�Pt&§g�YF��H�査½ƥw�s8��w�t�ՠH�p��,f�h��`|�(G�>/6��p@�����ޒ=hu��G�������ֈ���Ѵb|o�ē��*ImBI<�;����5�	$'Gе��U���[�E"ͥgX�1��&�eC���<ɇ�k�'����zɄ��r�7�pH�%�;�~�b��H�~��-�1<g��L�5�����#�G�D��c%#�}��N��� +�3~d~}�ovgA�W�~2�⼼����v�!~2�)��T��||�K̜���$�%�+r���·�PɞݒJ�O$9��|����sZ�>�m��	D͌�Vd�e��$OfD)��!��$�v-�Qd��\-�e`Ѽo���|S�'��"���d�N�9����b���Du\�ӂ�����+�;�{;Qޙc-�,[�X&
ZΨ�NqQ���0�"�'-����5��+1��������V��q��$A7�B����=1p�j��v���xʋ�(�҈	�����!�&:i'츷{%'�\�&�[X^-��L)���l�My$u%�3xc�'��>���J��5h#0g�
U~��0��䌴kk�hU���|[�̜�؃�	�Ȁ?���Ͼ�V ��Eg��C�Y@}"�iZ+eD�n6a�[�2NFs�4��_g�� 4��P2�s2����߼�0�2@k� ��.D^�s���t�(娕#=c,k�[���ޒ�Ȣ�Y��ۡl�R��m���r�kvJ6�b%�)�sGy/I�M����o=6�թV�&�p�+]@��'|�[���^�c�L�;��-M)�[pM��J�VJ��Z�Y77���&���� s��0*K$�!Lj`�.wHިo�ݖ:E���ǜq��sl��~b�۪��(�����IDPj&3�+:�Ιì�����Ae�_�_�C��i��#�Y�-~ɎL���[�Uےn�0�RZ�2��]fv����x��BŃ�֒��0ENpR��{�d.�:n�G�6F��4���]_��-�/2H�6Ϊ���_�����+&#k#�!Acl��/��Ku��'�F�Q�Şϱ�k��<�
T�]#|�+܀i [sr��>,��\�I��.N��Tߡ��W?�txvԈ���>? �����r�}��Ʃ���+1$l���6w_���;�