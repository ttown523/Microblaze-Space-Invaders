XlxV64EB    fa00    2b307������g�������Z���_�j����A�"��eq��y�Y�G6��ǩ�jEs�k��~��N���)���$93ao�|�ˉ9�j�?�T{ބGCQ�c�ST��_h��������۝ZA;��9T���3�/8]�a�6����$��Rz&���^�Nn����:����ߥTe���-FaOS�*��6�֕\�����"/#��[v��`9&$'���V\Q����Hֻlk�̎ot9�Ȟ�#��"C�\���Z4���fkZ?����h&����d�c��R����S/�.r	�1�=���>�ъg1��x�s~qu��hS
�P�{�����|������gߪr*�"֕:���1't\�#:����\��T�U�4,�]��/�M�o-jLb�e�w��)�*fhp�jA��77t Az58~�}~�y?�ɖ����_9��qp{�6#���(�ԅ� �~F8X�^qD˘����Y�Q0�ݙ	�ɔ��N?��0{�Mu1��P�:�f��|��Ki�X��;	�����N9���v���I�+������3�"e�mk2�J��zj;�����ɱ�̫V�5���qқ4�������I�d0),��||E[b���?����s�y��xjg'	��/�*�Ip��������]h�!�E�'+>.>�H��D��՟��	YD���P�|��i�w�;gpY�Wl3P}'b�B5K�C2��K#̧)�Mҙ��q��	����0�O��T0�	8�k��I��4���R���嚴�T�iQtT�g)w�>�n$Z�/]Fȼ^@�{1�O�`�z^��.k�9�N���@v��w��%�u��Z����+pk,ݑ��k�N�	�f���_ϖ|���(�?�?�OO�fuEt����(a�e���%Oz� o½��������D����2�9�h�E3��&��?�T�u�0�=�*ύ͸t��B��H\=�qd�Q��n��~������%��o��P��ϼ�y�T���}n��{���t��8��o{$��ۣM�:��X�x���P���)}�Q�iD���d'"f9h�:%Z��wT.}��&}$p�G�I��ت,�=��F�,��+��h�ۙ�+#�0���*P���p�Q@�f%�[_��r�c�^���L ��wi����G��g��& �5���B�h���̶��BJ��sJ¯	!"���p�
��B�EQ	np�
�Eƿ7)��\���l�
�]!Hx7~epo�
�p�p�EM1�/��9�SǪ�����[���C�t�
�?#: ��lG����E�gYQ' �*Ú���#��G���^�-����\�s�RE��̶��@��s[~A�6�'�BH���?U�ӗ�R�$���Hk���b>��}�x�#}?�uN��X�nfU��©�^��.����?�(S���X!-�d�DН������Ez���.���RPƄ`po&���]J�į�9���}��1s���?�_a�i��;��'���+|b�}����XUJ���2��yBX�ٶq����,!��\4cf�=�/I�V7F�O4E	΋�3�4V��S2s���������c|z���]���8@ٯ��)�˰���[��L�5pG�ڃ:/QYR��!��HU7E)�UEQ1��2Jz6�E���?�%�t�S�F�F�߾aߎ-k�Ǒ�7�W�S%Q�(jaM�E�,C�8B��+@�M8ԇ���5�EW=��Kuۜ�9�l����W�Ca�����T��e���*�u�r�c1��\/8"1Na-TY��}����p�{L�u]�Iu~�ЂH�����.>���c!H�����&)"l�}ϊ���܋�L^�����Xl1z�>���3��0�S�5����k��=I��B�l�-�a�`�\ xzI��i���@g݉c��6�#a����4ؿbr�1��������?b����xx^�o��iaR�G�0n�%_��2
�*���)�g�c�}�} B@k��p��q�1��ɩ��M�d��L*Zy�*����ڗ�6�-�8֤E�"�2V����Qk��Z+�O���["Y-:�䯅ٱ�a�1�:�s���[�f�791$��J�맍�h�k_�	��'Dj��{�n������3�i��6"B�j,ج�DQ��뷾i��c��_�t��c4��α[V},v����WV�T:��;Xk2i���J��n�!=�[N��T��w�?F��?b�؆�+n� T�]T.5-�N0�s�l�?����֤��v�m��ƙ͵��c��;*"w٦�,j�@��v�v����x'1B�u-M����zw��x0�dX��ڴ7�Ab����s��x�M?"���݋���1+��_�2�3�Cy݆�tC0�c#L�� �TeO�"��UŦ����:z%�g�i�`�駘��Ǳ�xƽ5^O	�ߐ�Y� x�}�t�ߩ��*6�h��,&��U{��_�K� a%	y���;����W�`.p���2��*yn�]����ܔ+�����ܫu�_�4��f�����9�=D��g�T��+W]���[5K*�דͷ6T�6KS��!�>�a
�}�~9�i������+-p:Oe����@�1M��[A�U�O�������"�[�)��,v8[�����-�,�Ѭm_I}�-�T�̸�+US�d84,�����Z��Ŏ*E�"�6U��@E���/��3=1�	V�5i�|�����e"��i�)/$Hpr�ʮ7��}�	c���(ה�d����p� �g3��&�����#c4�f���'�k����O�Z�:������6��ts�S�d0T�	9:����G��k�K^�#'.Cd���1`T?�ͶeS\3'�u���^�A5���l*Xc�&��X�ճɈ��*5�Q��Z���ܤ����o�}�CzP{jbuN�lvu	�!��*L��Ъ��QvP9� Ң
�jŤ;hn�"bn5g�".�:�+�97kט6�϶���<(F�}[�\Z�&���n���wLf_1�^����4i ���3OΟ�y;�5 w"�^�V8�J2z����b�..�e���#�Ÿ�p���P+�#x��/�X��-,5�e��	%f.��F�$��f��V����H��b�yS֠�A]_�aTE䲰�oXڇaM����{h%4���9?�?<d �lZ$n��@:�J���e������.:Q�
�9��um�~Z>�ӫA�2�wc�{���:����,����K�ȑ�+��ʰz>��Z����;����٪5Z�DF���G�]W�8��z-�mC%�X�d=Yŉ0H;t�?@�,Y��{�TwX?"pC�O�D�M8ۯQ��ˡ$9گ�fhM}cR�c�5���x��X�2�����E�6,�����'��� ��O2UQ�������]ـ������b6]�4isG�W�����קɌ�� <$e�*a�p��Vq�<5��(�M�R��V��id�ڛ��D��  ��?�b��Z'�s�"�!h�Xѩ �ٍ>;ON���$B�%x7>���EUF��{2�_�%E/�����|\S�ŋ�#9���En:�6EL���sʵ������)	fpy'���@�{I{k�N�nM!L���7��O��7bd�*0��U&h �TJ���x2B$���;�u��,U�gA�"	!���y��� �f�p'ɳ�#�~>l_��ٜ�cJ�-��]v.���!M��q��P���A�VP�� іZؓ�bM0�9Ϲ/��hQV��b6Vj����3�y똤F�����/mƑ$%�"_{���1���z�������� �P�cT�!`Q��dwS(�sZ��J�/���"��.c�!ج�^NW�h�y����9X�dn�#1��6� �b�Ԛ�(R�C��#�j�M����^�����(����޹�/�U+��s�����m�5[�q��[Y�k�����V���2=���ڸGF"�~��R�0
ډ�����T
��Tw&!�K���֒�&'����햟4��a 0���6�;~��\s=5����\��ӕs�}PZI�����ݤ���Dd����H$Bֱ�-=ޛ$k4��̺�:̖D��q�������3�B�>%{`N��$ �5`Y�����~>�'�Ɵ13R�����2��)�����U�ޚĂ`DĂ�H��~�2v}{6���0�-9�����CH��)�b,�RJ� %��ͯ��(L��fF�Ɖ@Ԙ;MjL~K��(�a�GSΠ����K�ʪk-�*r8�=#s��6<C����O5j��f*."�x�����p�Ce�~�"*��*A��\p�+�LF�0�͔��*@ɤ�W�D�hS�eB9?��Lh/q�Z�`��^\v!�}�����򾝀�#��L��!k�Wk"��N���&�<�d�2����k���1�0����z�{Vx�<����#ݚ�M��o�	a��A����C���!��Hm�wpIK_<�@Mz]�N|Ѿ�Ѓ��NS�f@�.��+�Ы}k-��H��'_�Z&w���X��,��O.��f!��.�G�^�����?lD����'Z����������\�Jߟ�|-�̲!S^;<���̜]�]8ֱ.چK����L�b���D�mM`X���]��~_���Ց��K��б#��7�xI>h5�j�!��k��m���b �o���<1Q`�S�2�y6;z`C��ދ�7��lAL��U�"lY�):�׌�������a5F4W�({ bX��@��ֳ|��4�}���?�q�.�v�V@�A�)mɽ�Q-A�:�r��eAx-;�s.�K���~��S��n@�9W�Fq(������j��'�����fZ��2&�|Љy��EŁ��CM�`y�7���\~IQ�$X�Q(�!�lIP�(�AJ�N͐c�]�~���o���� :(����H>��W��UO�ٲ��H����Q�`���b�2u��P�&������3ۓ%#�;* �o�g2����Rs�}�uK�`�O��戛���
�n�4}TĕZh;1�.���s6����cJMmj���MSC��|#�CR�����.�Җ��.�5p��/��vݦ��z����R{^s�.�N��f/��е�QS��,����[����XS����vg���*vj���Z���%M�ʹ��U"4gz:�� �|Xǿ�_�=/�$}���r��!"�!��y�D��k��~�\߳\�X�韵45-����5z�%~���ڧO�����U/��B�{Z56���n�X&���ۅ����+��Z�ބ�?˝)�q�*�����cO]���"l��K{�����p�����;}Ȭ�e����t{ݪ�ʝ���B}��D߿�G���ʭ��ZG��M�נ��_�����i�[�~�e�]�'���T�]�����լKIys	����'�v;P$?4Xgd!{#�@������,e�1���F;@�ݺp�+�e���%!)��u.	0"/�}��j���aGP�#��k��5B�2J��WqT~$��@�LJ.��N���rn{^4?W��OM��x�~	�Y�W��`Y�[�cc4l�"�%�.of��^�H�r�&���M�i�6i�ȳ1^
\R)�&2q��\�g��֤���z��D@���O$���£��.h "I�2��YNa���*���8��
��LХ�;X}`�� ��0G+6P�Л ��5������2LG����2'��>?p����?"�]�c:G0kV��a���̡��Ϊ���i������$�%#z����=���F?V['�=/rng��.��K�
b?�$bؼm\��t��pS���y�T#�ԕ�O0Q�/�y�S�'K�*�Y[��OȤֿÔ,�4c��mOl9��]�����=�%�Џ|��}�A��Ova�l�k����F��Z����z'��Ɵ�nUFNp�
$��C3���,tvKǑ��˘孛�Ʋ��cO��9��m�8����d�T�O;9x4�~^ƷE�)�u?�JR���A�K�� ��E��{X���0띇;�3όɕ�鲟�@�ې�7�gK1�7��7��^�f)p�M���$B�����A��F<���A�╅ x�3ڙܝ�v-�k͕�=����:���N����1H�)�9DO<n���taJ0�ޓ��l�fDeq��q�IhE��@�2O�A�Y�Mљ
lޥQ(&ӑ�M6#p��i�V|�&���K������&�~���LY6�� �C����t��;QF���A�<Ȩ_Fi$���@\���$ʢ�q��HY��׈(6P�=�cH�YdO�~ޑ	;����'��hw ��U;�LgZ�D	��*~�X��Q�Ii������p;����8�w���_�N�����Ɇ����$�V�C�\/S�	�%<	Mvs>����17g�mR� 4�۽�J=��n��R�уS�!��^�Q���Ŏ���S�Z��M�'B���>����t�0�0�� el����X��ъ�(X�ꓗy;@*�g>��j&�΄RaϦ9�k�%��*`hU�?�!�E����i�=?Ei3��79��)�_���ie1�R�Z|��ECE*�ֲ!�|GAMK��i�J@��{�;-
��!5S�|$s��&�ʹ��k���cp��%Yq���{>�W���ޝ�yo-[�t��>�����&�������e���=a]�d�o�SMdH�K��Ίu���ݰ�䥏(#�0�Bct�ቪɃ@@>������i�<���CiS\�_��V^����Zb�"7��IBI-
�lO[H5;7���u|�̀q�T-�Ok��ў*�@b�~�r�T��\��L
�&G<ԟu����^��|���^����k83I^Ǧ��	&�#VU�h�B���08�2P����Qaa�
���k昁�!�.ܱ���3x��[��jb�$l�p���
2�}�{��w�pԗ�ݓ������\w��;ĚV��:�x������������^��!� H��{�m�1hE�G�ޔ>o�خS3�1����k͏�G
KJ�]%�Ⲧۿok��fNWІ�%s8�`Ԥ(�bB<���F�8�nS���;�NT�@ "T���q�c�����~m��]�<��7�(���Q����ݸ������.�o�.�55�+�x�<4���eIh�#M�z5�4T�J&��GK��Y�E7o��܁C����C��a�|�sh�-.�![�{t[�d��9�ۂ�njv��ڠ�j&�m�R�7*��B�Gq����Ӵ�E���O�%�:��&��!q���ua�Q��.;�Ҝ�R,��uj���5������}�J+

� �?��/���P�r�,��k&���t�B�����4���đ�Z��M@�߫E�V����1����%�L�!��� ��v��)�n�H�26�/��G�0{��" ���&$�G��oo�+\�ڪ�d'>y**��V�<�T�ܿ�Y�8�Vx�������&�����K *�D�v*��iQ�q�m�}>mY軩n߿�1n��)�vջ3�&��])�(7B�?�� G�V�M"���*	��}u��L��K�ﺒ[ۡy#+��ǩ0��0-�F*_B7G�v�7S:ɷ����R��� ��ܡqF�j�a�����n¬�`T�]��;�^n��[�A���^S���8��4&�q�Y
B�K�H�Iu��f`B@��q�[�-C���H7_"_�(���J���%���~_*���������"���D�;��D^�('kr�^d�)��7U�<�X@r
��"��Kq<��.�P�P��#��[�(�������5mw{
��g���v�k#�!��T��^��t��fJ`%�lOKǆ�v��O�(�K�@A&V�%�1��A�"�|�Ֆ�8 �#LO�/��<�b\�@&ClI����E-37X&i^M���>GE�����&�f��C�YO�e���?Bw;�HY�Aܧ���G� ��m�"�!~օt8��tF�6hp8q��uuA/3�dq�+���VD\0=�g-C�C0��pPi�-�
30�77�r��ݶ�
r����P�|N���ZGHK�^ԸV9S���I���=�+R*T�����a+���A��+��zR(���I�TP
,�i_�搄u=Z��
���+I╅�]���ON5��O��;[9w��!F�=r[wK�����Ô	�_�����?�sF�NkZ)*�LZch��b� �\�����ճV�R+"xL+|�IP�K*�)3�x2�W�|�C�$�TI"q���a��	����:�G�&PyA�䷇$y��%�f���厪;֜t0<,VT�z�В�;�87'�Ht��N(�C�o��� #�e>΂���#�cUc����Ygl�Ԃ\	��b��������`lY�W������/�m�a�H3�Ǵ����e��q�"\�}te����j![PLJ)���,G�?Yw��7p�<0wR�!/b
�q7>ώg���Zt�sW�л�nSE9���U.ㅻ���K�5C�Ś�|ٞ0Ei���
��K�o���?�P�[�|�g��#m�.�P�ksA��&'R�B��lS���d�7
=v�3� `56� �"���@i	��8�QH@7I�����P�=�������{��e��v�G���֠�=&t����>:fݳ���NJ������f�4@䘲�'��Hx�Y�gg�+v�b`�d������,4A�gia �p��d���B5X�:��P
�T����+ׅ&C�j`޳pm���I<.�'-t"s��ڍ�1�7Yj�93kƪ駂�����9�=b�?�c��#��v�U�$(�֮�v��n���=l&F�f���Ǔ�]�`�k�8�hYmu���s��Hv���?�ܒ	ǻč�O%>�\w� (��f�ᮏ�.|zp-<�;�w�q#/t(g�����ls[��Pc63r�v�-�@�r�h�P8�$=v%��x�A�{��A4��OX��Qy�4�rSz>��d�ߏ*\���r31���x+��ʊ��	"����O[�������n�0�x�d*�Xɻ����D��x�n�K�����e]���9�À\��*OU��X���$Ѧ����Z�r�H� �LΎ�ofzn�	�#o%�HX�9��N����|M��Ȓ4$?������$	��b�|�g{�� ���A�yP q5����_p��#;��^���=�k�W���A�G���aN�Z��u��T\�ر]��39��=�G�;Y)%���H�mXE�<��-n/k�Ȧ�3|�<u�OZHG�ai�
N3�g��_�=�7�-M�O���
����B9�v>��j�2�d-�h٘Sޢ��κӈ'	��	�;��r9uĨ�"L�.�PK��AWP��Dj��rI\�������Ε��̉���B=��|2Y$:2���W��t���c!��N���#3�����dm�8	e�;��_��'S�"I�j)��6	I�$q+����+�g�Ե�,��]lr��5�)�( ��Y��E�a�k�z�Ec;�^l�"���oY�X}�M㠩�6:��m��!#-��	j�5�~ø}/Vb	u��t[-�Jj�K�{�7I��w����(�0×0.��EM#B�\.Ѹ�\���Y��K(ｩ��n'Wd?�(��x-`�!�`"x��6l-A�N����L������0���ڢ��^� �-�*BB$��oÖd���W3� G%\Ia(D�$�Ԓ֯��*g@6�-gɜ}��q�!�.v�����h�z����6d�|�`��Ă�ͷ�ؿwmp������Ԁ<S�1��6| ��G���Î��F)O��!쬸�y�� �č;�����c�����>�yB.��_5ՄO��_\/���}2��~q�U��K��Ő.Im��66a�����*��BBtm�y�u��gz��$<�#���v��`|�O-p�>lt�V(L�x�9b��;puX��U���k������k�C�aƯ��YcA��cQƦK�`��ݎxL����!Ӟ�}�ʢ.�d��"!p ����WQ�\�l3� T6��$�?�
��6�@b�j�3�sAu=c��6�(�IsV�Y��B��5ZQ-���H����s:p�ۨ�8��>�D)(`H��_Y�
w�)�Z��Z��mj�K�{>� �ް���B̂c!Q0�k��Q�b����3�d�E��1��������}=��J�Hܧ����6L���mo�	ɼr�-����j���9�Y�T��F��卤�_�#�e�����_j���?�X�>�qH&*��F�g��sYg�^�q%��vk"1D�f��D��P/V�,�k��u����m���j�$6�T����s���=�WCOʷoIf�RmA�C:oG�9��l���%������ZZ�m�������5[&BUC��-j�����NE�� 7X�o����o�b�3j���D��L�ɉ���Kh��C\WM	�V+ԓ��(<�l�炷1�ԁu�/�W�a�s\�0q�I����6�����H��wOk�Ś��p;+H���ӱ΁�j�|kr\���eJh�*�����@Ɍ$�Ŝ�o�4���=�eW�����^u�l�N��'Ϟ`��!��ȯ�MlBJV�W�Sb�����Z�j�L��'i�9�U�i:��*�h��X�����Ҥ���V�����ű���ϔ��Sb��\��؎��Q�C��\ٰ�޲���L�ޟ1��T�M�kH��4\<=~5BQ���*��N5���v;�87��+�{�"�NH���i����_?��|�1U�9����v5i7EJ������<�j�����$�g�`҈	XlxV64EB    b8de    1f00B����Qڈ5�� ��۰��s�E�J7E �YB����Ɖ���>��[[nv��۹�C�L���w�l	GC�*�a� �� F�!��X�Q"�0-�R3:g)E��¢	��P�6�i�����}�~�rU���D�Ç.<�-�Y��6&��1��[�UNp�&�Y�?�'�%z85�&�#�8ِ�P9.��#���fؼݦČ�@�+�[o��8��H����ܞ�;i�@��U+�r�ƿO��(��>��Ƕk^���w�2y�ǚ5޹HN@)����j�j6L�%1P ��� ��c0K>Vgo�ޑ*�Y�/�h�@|�k;x}l�&2�\jq:5����鏪3��хm���w4�4��A�$9�Ҋ�!/j)5$���I�/�p���.ձc@�������%EJL�Ԗ��{h`-_O�v��j��
�6u�2��>�T",��:3����y��M(���sj��u���	p�]/%�V��VN>{�qb������W�J^�rT��o�G{��R����G!�/z���������\v��V��,�ބW2����J��*��;ن�&+��R#�e�7o"�c?�{�新�}~)IJ�6$d���7*�8���ֺ��)��y�_���Q���tJW;�Wjk�z �<���u3�%9����)�A�����ʋw�F��ָ\34CH�R|V(��<����`�I��i��P�C	 A7U�s���~w�؈�p�st�R���@�����u�@���4�@�T�0��f�������/..��D�tQϚ�#�]S`2��s�C`�j���y�Sgyw��+u6����Q�ɲ�mw��qKc
ڍ�&�Fs�����|�:���P�k�J��KH�؞��;������$6$~�s�6kkUW�@Q�J8������$�����D�T��>$�*�54|�qK�藖�.x9����0ix��gn3H���!F��R1G���R�u�Z=- �g4X 
c?�W���:�d���i�F���R�B�����".N4�Qb�Ezv-�Bp��(4�n�B�!�e���� :�6��y9���czR���0nY��#U���i�ϓ��`�JW���z4�Km"�j�!X�ą�J���w���<�yHcH��@d�+��,�Iq-5X�;���צ�7ͳ�:�9eT̃�@��Դ�� {I��I��}�̱����1����P� E��e�] ��G�� e�z���ߠ��������zV�l�~�5�A`��SGM��{A3-U]�8lm����AMS@K�����!���J��\�#�'1}>�	d��p��QQ2mv3��+:��Q�.��[G^�>�Z��r4��2����h�1흥L�$h�u��u�ے��~Gf����r6)"��C�f�x���-)|�B-X��e$����;���/�� �0�#�o����!������N�3z}6�.�ˇ:��a�pi��X(x�Ɍ�e��i{ǎ귣s�ya5%V�n,}B��ZF�'��)�z�}/�[1O��A��1����4��Cm��K�?b�)�ô�?�/�4��*%�\��M��!}��YL��Ղ�PTڛ�eI0���ʯ��g�Ɵ*��U*/�uo����f�s��)�*M�Z��C*�� �Q��2�A9�K�>Z�����j~F����n�����iX��D7�	��;]�N�~I���c)6Y>�q��$�J���^VmH�ny��yω�[��lXLjxs3��"Hމ�xi�#St���6H��d!��9��?�Ѭ�% f�gO��~�fŴߊuppf�H]~�B���d_�ꪼ����j��P�q�6F��+�;Wr�Gl�Ӎ����̿��* ���f$���q�H� �_q�nE��6�)��טs�Mb{�T�n0���Pd�� ��0��v�w����	���Bl��]6D�������_o#��,�p�sUU%9�U�h�"�"S�yv����h�ZQ�ϼX
���n�����N[�V���/���>����UAP�/���\ވ�С�`�RP�#�|���5Ze[3��SC	�>�Kr��а��t>,���~i4��)R���NqT��7}�{��]m��&"��7��.�L�Pk���b�[=I��b�bg�1���4�å%X�f�/����e�()H��D�wɽ�w�0)8,K?Q-񑂩����ZT�˙gy>l��{���`�0�`�cw�),M�������	���/�QzT6)R��R7���������Xx[�u�π�2�ķ��j	�x���J(&!v#�Q�)��@�Z�^jqIiu�g�	�OX;bN'�\K��x�u�q@? lfܲ��h�͝),���p��/x�c�] I�݆������{�wU�Յ�r�.�~������*��r]u��&���RHP��ǫ��y�zj
d�����P@��E�W����bw͐B����e[��Hy泳��^��!����/	�#��<v�UȺ<%���V	4�T�zg�SV�f ����)�f�4��<�-d�����n�GR2%���0���; Zm��R,�_*��Y9��Ǡ�H)�H$IFa�!8"�ߒUs�$�2��m��W���=�%�s�2=��L��M�mUKk
����G��O�/��\vGm0�|#k�\��څ�A0�޴T�e�*�����z|-M�A�i��91%��8:�w1��i�X�llq|�m��3 ���M��b�~��$Us��B�dLg(��]�C�(�^.�k�L�D��R� ��I�k��h9=���F(8�:h���X6 �T���9}WYjːջ޳H�Y|r�)��؀d�M�G���_���#��ى�
9v����\�.Z!Ja���� \�;�8EW�*Ç��H���ot�5��\k����i��r
����R6,t.�1��Ń��'�9e�d��w����y�S[Ō�����O��MH3��L\�(��B�y/���$:�Q78�v,InD<�f&M�r�����{���s�	O��a��g�%P~XOWJ[�U����*Vb�]ʎiw.����ψAcY�1��+�
UDFE�w�6�]�`�[`�����Q���L��aw�j0�4	D��	HF�,
v���T��1t/����猎�>J��� ��/�'�e��=�3�ĸ8f��Q����Y�rd �xx�pAj��dt��(��/�����l4���ɱ�nR����2�#�q�����4��d�������$�=���Ӆ���H�=R����'JJ� �C�U&��|a *d�I�۞���"�-B���s�*g�N���0%�*�
'{3���$z�+�C���u U!��u�N1-$5��TP���:��6��DI���Rm��U/լ�m��cl���d��{��G���!�E;ul]m�UY2�q����r'�1����y��iȣ�uTz��qө6�b��[��`��fWY�çg��������^S���8 ��b펇7������>2��g�7h�-�� �^^yt���(G��^G��A��_�?���.DO`�wS���g?�ǆ߫���m02���ڼ �N@A��[�(˯�O���y��*1\W�zkA�Zd���"�O�꾄���=���c��6,q���Q$�H탕���o�ʎngh|f�'A�g{_ֻ���9T��"��}L� J�d�������OC�CjgaNq�<R��;+��YRF[i�� ��B!,y	���jN]'�\E��rH|
}�o�R'�3l��9��P��i�Q�&M�D��s���[\T"�SyeX�`�l9�<�Ҕ�M��	��*��������N�|[Y�NW��ݝ1&�qAH�H���;/�:�+�V
�E�N�h�L�KF�+�������V�S�:�KNo�J.���΋'�� �8��p��#^.���Q	� ����J	��r=����͢S�U���[<p�im��i݄�f��w��Y��Pt�< ��_�?�BU�l��Ǫ�u�\&r��I]�#�G�J��	`{�Y�~)���Hȋ��X�*fj����s�îx�]"��-�i�u��$���9��l(FX^cԂ�@�p�qB�-~�$��An8�������`����Q�e�dm�C)"��P�V�'�Dan,U��DVp�����mdWŘxyFN�c���O����q�ַx��8����3	��l7FL��T.��K7�v��;�&J��͗Sm�q�&�7��a{\H�m��3#fIh�)�V�ڋJH|�2�zO<�O>|�m��{���ȴ�$�p�$�p�7�uX��ԭ�J�k@_eL��sZ�W�i��RC��
h���)�!:���J���̽��a���t�%X�)R�5�Ŵ�\��ǡr�M���a�"��$f�:1�XQ �4�1NӜ���,�&�*S����JҢ�Kxms֭	_Olq��'����v��V)���ᘷ\蘠�2eV���W�L)da�Hp8G/vޕ�θ�n߽b�|Wī͑�cH��B;q�{�iu�Y���<�cY����G}/8"����;d�3�I�֊B�s�éGU����6�3���h�7���*�Ab��dPV��:8�&�O�;�����?46��A����YɅ*�PR{yMuX�K�f�4Z�]���] YP���.%i�-d�Dւ� Sn�n5[c�nK��=�`�4�U���"��?ބ`�Gٺ�/ۿF�|.;3\��l7�	�L>������?����6��hߦ�/֧���G����t<Rn��)�;_�CVA��5d�u2ТAb�����!@�e��RA��d	�آy��HM�ҿ1�o�3����ܷ�4�	����Bj��c�_�)��$��*&pX�i�aK��@��m[�$�h�)`�FӿI��?�ේh������@G���Q�Q!�0�����F�Ai�0GfNf�!	��p%[8BǴ2G��S�I�$��e��gO/�JN���L-����-E�����ER���~ڳ�F�$�%�eZ�<yR�G�������7w�;z�+�H �_�g.�n���R����A���6��%�:~��
�j,�c����k'J%�D	
��%uN�L}��wIC��-�����C�lP��|�U�q;����W!zy��z��U4+~�>c
���?H�wc�4ƥ�����Ȕ�C��e�&�)���X`�������/]N%��-WT������!!���Y�G-ML�r�YN�]��s��A$�D�v~#G��/V�b!
@��֧���I {���L�o���^���v�P����C��ҧ�E���'�C���X�k}t�c��T�آ�������9�y�Y��ȍ��=������#a�H��#DK������xxŖ�zE(��e�|k%\0���l��lc�u��v�dI���BE�};��W�6@$G���O�LLR-�"�!�;�"����<���T��R� 2�{����*�+t�5#�3[�:���(��|:��'~�_��r�%�Ǟ��FJ��u�!���w��~.��̢�UL��J�gz�@��T��Hi�����i
�� ��� '�_��3�����QLi$*��<�)]@�q���K����8TY��"-��VWrU�Y�W7���\�8��!�]פС@���ߧ/��1^9���ߊޮ'5T�IIzV�|���y���覱~���-�����0j����_�a}o; 2�7�F�AS�j�<^TИ��a�~�
�R� �ݾ�hd}SA�Ɋ�\E2�Cj��w�+�}V�5���B��h5��&5���4���՘�ݿHA��§ Lty�7G��86Z�i�Iv��7 �Eu6�]ƚR����{�aX�j�J��hh�<,��B�7ȇ�`5҄��L�oX������w��+g��&8q�
tk*��:4���KB��F��X9n\Y��v��w�5u7��$��C����n��}�����`S��^��"_膃 %�7�n��5y�PK���3нxWj{��=!�򘥢�8�J�P�H�e��:�=�^i.��R����1����N&"[�D�����s4���/�ψY^w��H�J�~�6n:�ӌD��kel.�uʰ�s"q�T�M�,{Z8U�H�h��l��U�╪x�WJ8O�-��%|u��$�M���I\7f��[;�1I}0�)��̺wE�2r���o��h���onY�,A(� �L���� h�J�)'��U4�-<:�ܣ�+E�6�NY�(#��Пd�x��t� ���s��Z����ǧ�����l���c�J���fn#����nH�
a�6d[|��\&��	����9>Dy� ���>!H^�o2�POr���2P.�Z7�F���ɞ�,2�GCHr�I$��~��n����:_{��*�yKB�.�_��qfmcN��5xG<���;/ϔ�+�b��B�d���"�9��3�~A�x"Ylu\\�K`�L��Hбr|�׹	^q1^��0���USk�j��wt 1���6a�ő*�G+�|��P �Y�>��a	<uA�����K>��K�^w�?�o8ey���ə��hh`��5��p���W��\�J:��g���J�%��
m��p#�%!"+�%'��:����}�
�ޠ���`6��fՠ�gP<��	nS�iڱ� �xm����u��4��Y=}l�Y^N�@x�23'q����sY���L���[�D����J����9`���ebWi�����?�d`M�����^�:�a���e""vvC�r��շ���B�5(*QG'�1m��O	F�(#���t�=�%�;̪4*v#�d���̙Û�\��66r]v�\]��q]aCT�;L
���]H:^j���gջاw�v���=�#4���=$!�mȨ}��� �#q�����@�'�3L	�j���U���]���SB��ch����CgA��[D ��]ʃg�i�Od�@�vj(i~/���F�q�iD� f���\u[Y�����H�"��R.�^�����}b����;U	������$�?�I"���oz�99[wTF��m�{";�8��{�'� l󶒉�B�芜e�FR�I	Bl���ļ�����T�n �a8��֢M4�V=�R,7��aq_��@��QS�d'
��$��2�`�ؤ[pʶv������߮����-��yL��/	R�����P#�؃�nF|�o:P(s��9NZ�N�����f�R�X�sQ.�3�)��y�����A�Uvܢ┙�G޸�lk/pq]Ǽ�KX�SDC�F`q����_���.��E�{Bu�`n�dx���`P���S�����}l�r��8���Tެh�������z����
5�j�S�
�e�	F�H�3'e����ۃ�B��^T Ny��
����5���,�����5˃�������h��v�k��1�N-h\�([cFDC��+B�6�m���Z����*H�!��(����(����K���R׵8��1��;Z���nOf?Y�XFi�
�3!��wdrq��~_�B}]� �u��	�������~��(j»}��*!̮�O?���c��8@�>�;lZ.��7�tDP�V�ws����^���p���I���(`�,p��m��[PT}�qD:�	w-��}�)g(�2����Ba�v͍��,#xA;�i ��3�>�~���P��'�_�����?)