XlxV64EB    1d2a     9f0h�V湼�~��q��He�|�n�w����hD���~�z��;� ��\��T{1�2ݏ|�c����1�����lI�lQ{��۹X�o��w��a��o�ɜ�91}�2�G!�@�'.�\��
��rh���Lpݖ��G�1�d5�̓aQ��r�O����~�dg=a��;Q��ɇSv^�U����A�`���������g:]��2#E����HpcZ2���Q@��eo�$&�l��s
+��c���-����X~�����`d3�}BRe$��4��OT�ד
���mm�
�K3�kI��6*y��喼��A$#,�J�nf����V��pѯ�JV_"���^c�yʨ+B�u^��|��8&�z��!ĳ�I*_����q���\~՗O�XG����BIc���(���<iؘ��u\���L�(}x�������޲;	amJ}���N'��c$�x|�>D���B�,�Ob�U7����)U#=��  ˜�K��\u�\6�+�"��HmǷ���,E� �eM˱n���� P།%�h�����U��>��=F��u6,�tg��W���>pI[Q�b�`�Yh��Ҵ�7�D/�ҽ�;<��$�oq��_��B4͢�P�m��X�.eH���l[��1�BM�+�2��E��y��������!�}��8��9��]<����?ӈZ����A�!�4m!@�F1�
�v�ˉ�C4&4׫�l�����6#�m� f���k���}�J�5@�Tx�|�8��!����Php>�c�夏v��Jί"�����z�Ee�6B���RFy:`%�X;�4*-���4o|��b���=$O��rw��s�Ki^6�L���y��9T��HyC��ŻAOsҥvϭ�k�>��Ś�U*�:��6B�x_m��}�,Z�h��yȚ��%�[����m�5s��p)=c��7@F9,�3�� �%?&m�)��&�I2�tw�P�]Y�T綹��S �^Ԇ��f���F�[@�oRQ)Ӱ���G���=)�� %_��6�2�,�;�4�X
�W���w����}|��NseI
̣;�MU�;���d�;��_��|a;�p,�@�xpJc�qh�n������n�0l$��G=K/`'�}�����qν�8��JmS[c��۟�C�)vL�j�)Ÿ�:AG8<�7u���|���-������M�P7F�{��jECΝ�S�|@�����So�h"�oi�~o�x�}E�`�ܿ�gt�T���4}�0)����/����t���*�������Kg|n������X��Ze'��a���p^�tv��ژɓMv]���Y/�I��bsJr1�~~��I��(�9��d��L�ѺxY�[lȊ �ݵz;��9���^g|ُ��搠�D��ҩ�;�9���}��S(ʶ���$�VZ����bը���U p�4?���[�U΀�����% 6LB%
�
�V���/��Ce���HΆ	�6��`AK�&-۷�A�v����T3e�9�����Vc�2p����&�hvv@���H�v+(rH��䘵T�/�uj��=^��𥽸��&C�Я�AY	!_�n��*���&��Gf��{�$ɢB8����qZm�p�[�E��xG��-0f��C�F6����C�v�t:��&;:7��*ξ1`�W�E�nx�g�Y�NjQ9�����A%�>c��y��;c�f�>�ode\���]k�"5^������n��Ѥ/[1����C��um%��X{K�?��%0�����6�ɧ�S2�9������az�	a����;a�;���2ͣ(V5��H����*/�#���G�����~�b��?��m9���rj�b�������
�B��khM]���h/s��1��z2���S�;10���F��˃�S�����-Y�p��i`�.�a�9G��X��2�Ք�ar;���}�KYDRڱ"��@�s��i;���HaD��3}���ƆrV�L���x������eU�fuoYW��?�)|�d�E
�Fx�М2�X<Lh����>��>��7�3<����{�?{�E=��^�i�P� �{|�������"Ð'�,���W-34d���X#���v��wa�q.���f���x:}aǇ126�-��C]gfl�{�s��o��{?�k����^��[�iN���(��fӑD��t�{��C��-\#�'$�vC�=��˱�����9��x�(5ۗ�}�3CH���`��[�̧��v��Qa��f̧����|�xn�E�c�3+�!�lVO�`J��+O�&rlͰ�k������n�s������-Q ����vŁ5��'�!L��9c�]Ex��[���M��1����:�?�%�����y��<�)%�
#;`F��4���6�0o�z���2}��������[o2�+J�;�+��U�����