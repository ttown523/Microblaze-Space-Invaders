XlxV64EB    3203     de0�I�u�S Yw9���UFI�C�Y���I*pl7g�M;=g�5cE(�ب��o�W�?���f!אG8���Q�o:���%��B'
�G�ݔ8^���u �`��|��YOv<�7k�ozDs��wv7�8-SX#�2��.�Eq������);��%_G��Z�1�_�΅^r������!}t�pF�7�#��'C���[�����)g���T��v��o����&].�sɷ�]Z}b��1����&�~�a�3�-N�q\�tYJ��f���8@�;W��R��f`mT�Qd�9ӟ��y��]�J����L���o�
JtNP�_c�o���̭�䆯��Ƹ�'n�Q�`rƆ�?I��(�A�d���핐��ɮ��D�W�B+�|��&�~�z@b����o8���N�\rZh�x	_I���v�,̦�d��$F��Ï`.�M^�������Vi�����4K[��$��k\��]�;AQB`�!I�x���AY����>�!l��U	괣E�>�W̅�h�fchU^�t>WR��]S9:���0�ǚ�[��de��+�%���5
�R)ID�t��:s���2�{��0y�'6�´�B�as֠�hC� c"]��<1rjO�UM�p��qNfK���n��vS�S%�������}���QQ�U�lO��9��ʔ�ELk�N?c�/�1&@ x^DG�tɇ�wFtGSmuT�N�u�\;�pi��Lg��=1E�,���W�I���N8k ���j%u<�S�j9���OVi�$��?��D����rD=Nݤ�;;�~u�)�<�JN��a1����r��ɤ�o-�&�0�P+1<�
=���x�k��#s���d���H��/�T&�u��q].��w�o���+V�T;:�~���"N�"���~�l��?�2�͙��%<$z�oW���J,��Cڷ��=�!��:8��g�
�-�N�

��l`��̩�[��I��q��;q��Q#J��S&@2��hN��n��H_��6z���=�v�eUu�䴟���2�o,Pܾ�����$��3�*��S�P��@��D�p+���ï�B��论�ү��u��vI�Z�5�2D\=��o�fWP�����E��Y;��k֓�G��%kg�l�s��SO�y����)T����4ʓ3D�3 ]�k��h;�2��2�/p�"�Vu�B��3���.�v�F�87��e@|43웈��@���W�Y�m�9A\g�g�lߞ�.�5��cf	T�-��%k�Y���RWe�电Dʠ���=�/IT�JR���)B�MɦaO1���V�x3�PYEyz�HP�ڼ_o�A��y�pZ/����@�������'j����R����a)p�l��EJ����׀x���\_C�G��J�H <�!B�z��=���(o��
�H�<�*~�j;� L-H+�9���1�ӱH�)�5�{&��y+2:��y��d�/�4�*�;�+��&.ʅ�H|��]��Χ�ze��b#E����l����#���d�{��|��hV�~��J��v�/{Q��7���d�\]�v���4���ϓT�~�}�����Q|���9v�\Ԟ�P�0���<ᩑ�jQ��h�Q	�2f"�` ����՗�EU*SN$� �1���~::h�1ixJ!�m̽�+XX��U�@f"�,c#�\a��P G�l{��"��E�2�D�#�l�a�L*��:��}��N�q0���(�����p��ɕ(�߬V������r�%ɩ#7�~i�˞y-�$>�����|��T�1�8@��¥�#"%��:�Okp@7ލ�K{W���wdA��'�[�yƈ<]�1T͌1��6�V�� :�'c�#Z�Ңhb����8�2c٬�dH��ᛮ�jkǈ0s���.���ï�i�[�"\<�ݑ�@w��=�@_{۪�I  p7~N�2�1��-Q��Vb`^;ˌiq U.��7�Y��Zt�H�|3["���KB��mt�̙<�����75K+�|���JYI�◤��!��IG��hej�Pr1f�B�#�JU��w��3�P�Ot �b�>7�ڶ8.�V�EJ����8�;\;_��s㓆ڻGĖ9yڋ��܅z9:`Le�C��H���C�H��
�\�xAr��]<�_�D&��KF$c�Ea��"pA]@rsq*	�I�b^�5��р�]F����q�-"2qDxp�f2�j�ڟ�%u���ʻ�M�m!q��[���Y�y�z�x4M�hoX���Ne�i�h�*���{��>(KW��Y�.��$����k����+��e\@O}t�H�8CCY�'�T}������x���}w;��+����F������w��=��x����u!�T�ǥ>z�yjI֯�D�z��d��e��1�`���3�l�lư#�bd�g�=F�4XR����0,i�q�J'm�@B�FE3�Lӥ�A5����H�����TlE���?Z�:�\�{��f�ղ{L���{�T�X����v*[s�mp
��4a��o���1��bi���M*!+W�چ��TbVۈ�q�;�ގA/�m�O8�4��ֹqhIx�� G�Y�����T����k�4���B]St[T��؀��	�_����	��4���6^��W5��BQ�}


tAƲ�ҝb�lc�h����n]p�&��k#�'_O���͏Lns�.*��<0xY�T�S� s3�0��PGӼW)��x#۴^���C��>�A5�Y�T+v�����g���wX�{o��}/L�9���S �(�������D��e���С�}?po��]_�\!��~�yo���ٯy����4��&�J�����4������E�B��'���]����Jt~�+!G���#�h�=-�������̠������I�f*��(���=֯3���_�F�Ym��xH��6���t@�����,pal�7��l����2^��XQS��lu|7��pt.��P�y�7������_#��jy�!�� v��lfn�,��-�����TN�ǖ �-Vz�u��"Ss3Af̖\"}ᄰ�[H�Շ� k���q�]���Ņ��;Q0zhtH�]�,��?υ��y���s8�b�de���:��.\M�q�e��J������@a3��wX�?�\m�'м��s�ltly&{O�BE�(���E�r�w��S:-p����c
᚛��ZBF!�gX��\"�<y�Z_B��IOڀ��b�1�cb������c�"`���ֈi�����Dz�v;��U}���[�����,�ܩ�f�$*�H�X>�:�cB��t1��^��e�V��ǫ9T�3}p'Ė����{��ѝf
�9U�x,(>�mTt��_���xM^�3tkd�FG%?��'��Z�=����b�L
���Ǝ|�-����W��y�(M��O���zڅr����/֨O��kk��nM�s8w+'��p�0�X�8�