XlxV64EB    8b0e    1f50saf9����	���������b�[ĞH��J�B��L:n)�8��h�O0d�d��\x�D�F�0�f��y30[����BDÀL[1)f�+�TJ~�/#�\����z�vv���	&R�2�	r��Ď>}F�^��� !�܆��?7�V�A��#À�$u��qvP��|��~]���Tt�L�MQ�����^��HS�c�{��S.Z�K��b[� �u��&~Y|@2#`V�TƉ����N�p}�9�A�^v#��L��QQ�a�z0�WvP6&p��H�s�4j��n=����|H��D���2�*�C��B���㶌��$�]9a�3?f"Kç�[r�ޟ��S��
 ���"�)^�:�=����hh\�~P�T�Y�nt�"Zo��c���;%(}�;���Q�7O�*F��%k�Y(����f�At7�F����?�[�~
J2�d[�T1���ۗv8�O���ƹJ�6�P+U��شO�B�|M�<�9�)G���+���@��:�B���v�~;��L�bV���؟�0�gTs��b~,��OӍ�K+Sf���n�����C�1��"@C[�c�k�L��ַ�ۛ�y��l��`�7Hb0Բs~J.Av��^��k����u���)S���v��g���G��;��D>���\�C��¦V�> �	��9}�������OH@{�ɲ��/;����EՇ�Y�7�N$��N*�bX��F3��8���I`'�H��_%��{1@���%�Z�!X3%��))졗�βd.���,�ԇd�i��BD;����W��,�sk��4tC�5d쁖��J*tX�Q��LE+V��c�0�q���\��p�}���n�i@ٹZ*j.J?���Bg9�ϴy~��g�v���� ������d���}	��Hn?�߹j���t����K�,�/�͛��T2I"/R��7����~�I�B�vla�N`��ֲ�6¶��o[}N�d��C���?I�p��K�V֩(�G^1�ٯ���C�Y���Έ��;" -�8Zw�5��P�c�̈́š�j6��|O�lD�^���9[��꩛���FԀ4i�ƛ����1Zi^���]��:�Օ�75�2o�>��y�:��2)�uY��1���G��~�3,����*���e:��)�8�#-ٜêH�jh(!��z�����u�T�y�T��`�5(����(5O �i[�Q�ẖ�5����vW,��b�^���eЋ�jւ�`�
���GG�C6I&��?&��a�����'J���b��Q���VWr���p�s�wR�w7'�:Ĳ�{��Nuz}WZ���@\C�I����d�iZy�ŧE'���*)$~i@�l��I)8�s�^Q��t�ۀ�.����gFJ�}Kt��%XV>�rn`��Y�>�XiMs��^hU*�p��s0zʚ��s�>�FK�+���՚���d�9G��V֙^1�d�����@Kl,*��L����֜��^��;~�~4'GY̴�7�_I��<_���^;�?)�TZə$�
��o�[�kf�o�º�0u�	U��'*T!$Gg	��(��Ǳ�h D3V�pJ�݇۷��Md(vZ�����fDx9�,�p��3���o8�8�|!#E$�������rs�ؼy�-� {r�熚UhI�5�;�����Ĳ~m��K�I�.=X��C�|�����Z���5p<j���x�o���D��@9��T4����u	�JyEgX��0$�@���d_��������l�W�.��dlۡr�ݚk�9����1c��ip�(��������*h(ɪ¼T�r�(4m.�s�b$�֥u�Zi2���� ��ǡ��[��jiDPかIՌ.�Uyhe��?@���d�;��ȼ��}�X�T��Y��K`Sh�ԧh]�#<ț�缷����F�W�����"�����#���Ŭ������Φ����s+8$��Cń4�O�?����<��\�!�`�US<(�i�I�K��ݸW�T�M$��ES�:��
=;���lK����#�(���� k\f��<:�V)��G�߫AC�/l�L��veNͨ�s�]C����e�,&h�������� q�\aw��;��2~@w+|զ"	�C��h]2U}��{�s��x��9��n��NV�k	X5�?�z�9*��X�	'րP�ۯvAo�i�\�D<�S-�`��=cN���2c��`�%�d펯7	3-�W�
��U�o3.ԲkG����F+��?͹ݯ�h#a��,<B�.�!�!�-����[p_��v�i�V�Ţ�UN�OK�m�� 	����`���":rh-.�	����WuA�S^}֩_0h#b%�Ǒ��[!�#�����Ư;(�	B����M~�#�HzJ���(��{��y:�.���SO�\ ���{�>O݌_��!Mr�]찭�V8�Y ����ei6~]B�Ʒ鴹A5G[Q������[,��f�r�>�����j��k���]��4�|��������BP�Z9�c8�	A(�xf�yT����d�	=H�$�(�����#�=�f߲��$���r~KN����0���w�|
��`
y�kfE�=�]Hz.R�$�#���ѫ7�0�a���D����d\$������}�BW��c���?)�G�����z���a ~�R+�$E���(P��G
حץL�eU'�lF��d�Qp��j�1�D���L��~�2��B��q��ia�	sp�,���=�=q�lB�6 9�y���P�^���xtk���m�X}�w:�Jdr������D��$�tn��n=�k�,w _Rjѫr
��`s]Վ���������%N�׳6�B���E���`��	�7����N������1 ')ɓ�I��Eu������Hwl�������YU���>x$D��'�$��{B����٦'U�${ľ�eT�elٽO|��&�6��m1�y��f˱�J�4�9Ҩ.��~#��m���Rj�$[чz���{�l"�4��]]����.�?T�hw ��$��
�ذ�>:|?[�5Ư�-��4�^��:�Z"Gӂ��i��O�'��w?e�Br@�e�B���l��|\���|��!x�?/d]�q��yu�G�g�(��ƌ���I���UF�9,������2�}��50Q*	dӏ�S]͸4���?�/�B9�ҥ�=��y�U�2����r�Ȱ��LD�V���1A)� ��2�t!��wR��R{�Ig���k&�p1����(U4��K�"���I]�3@�Uo'�"�	�]K�,�W0�V��Qi����R���߲-��i�����.��ۛ�H/:��K� irK^�W�K�V������Jΐ���Q�,,��l�
���Zϱ������qs=md��%`*��D�G��m̞�De/�?b����" �����G�k��1g-��(}����۵�ٱ(��/��&��.\�V��w�<3�V��.��(�j?����r6.�0L~ss��x�O���{!h΂Ċ���\CyU@M���z�z}����Fw��N,�HM"N�[���N�Tb�� x�C'���1����O���<��1	�R�'a�ey���GY��r�Sߐd��2O+)�կb�����dv+R�L�Pjz5���Y�*��"�������8!�D����V<$1i�k:������e4A&`�Y�%p��	|����^�ҮSz'W/ �h���0�?3U�L]�gKJH���V% �J���rc���⽟��sm��|ef�8�FD��'������s,��L���}/�^<eg��)�L�J���@'q��T���4��f���Ēa�A(�G�4�@iV��Jq �E�I��<��-C_������p)9�+��3��1�娲���ՎB3 d��[P��� �&���jC.��o���/`V&�&5jlTF��M���AIbU����0��#���RD%S(�;���a�
ꋺ�b�E����5h�P���b�[�x��ug!�{L􆧮2,[��8������a��� �KB�pH����Vxu��xnT�ی�e���V���Sd�M��$�W�7�dix+%�k��{��J��~����72+5؀8EtYA�zAlc���c]�n�O�>���)�}+�E
�J�>d�9k�K���<J%�����
ut�Ѡ�4\��=�x��J�\�\�ǈ�,��?%�tg�����Y�~�6�9mo��O<�E��aaA6L��2If�����:@��$C���gP��M�4}�qL|��%U�p�FĜ��K��?�	��A�8�N= d�҅2
���==��cڬ$Q��9P�i�L�(���$E �����"�ҟT�=nB	�]�i�+�qw_�r`k9=��jaI��F^�r��G�r�L+!�2t $ťq��~+��{�DyKv.�nK!)ޞ�iX6Ǎ��0z��;�1n@Q�0�z;O�kbX7a[{�>Jh-�ɑ�^|�*D?�vmT�R��N&�f���������k���/��h:`�vP��	褆#ƫؠ�g�Aأ����y'ea6bͱ��{����c��OlD��44��U���S8����o�ٸ��@��Y�C��Cn�%��p�D 0� �T����vF��S��+�0:�N�Ol3j�h*�;C_P�@ P�	�0���
I�`��ޘR$Uk��ær:}|V@i�:
�A��mx��r�3�ŘVV&\�~6��M7�
�V&i�iD�{	�M��d5`��pPI����OUɷ�5^���g���D~6�27&�C�OW���/?�|�lF�D�z>s	6T���j����^,�F�������~C^�u������Q\��������{X#��2���TG���m��������Z�=#����̎g�l�}��w�ʻ�W�E�8#�I����~SpHb2)J+n�\�B��"_���T0y��֙#���%�V[s�K����҉W1��WB��Ƶ��j`.�����'�O�n�n�֊�?��(�$޹s�n����$��#e�[0�
�����)X\�Z���''�����c��Ifh�̎exE�i�b��'	�с�4ou+�D��)9�N�H���倐Uz+~*�5Bp7	a�AП��gz���'�?O�H'y`����N1 �p���X�NR���M�R��C~������-1��� �M~C�Fzl�Ϊ�Gt.�w��s]׈�ln��}aj��[k}����.�I���.>�N�LY\sB� %���5YY��I�p��z��cqXA��෼8�q)��;`����Z�nM���a�yխ�/�h�\z��(��<o�7�#�`��J�ł�xҋ8���t���d��ޫ��(�EkwjA�_���oG����(!��N|Μ�[QG�Xג���uKҚ5)���1F���z��D頒�F~<�����3f�֕C�0����p��}9�H���o\+� ����۸��<-�����}��Z<�e�N��3�2���ه�����M����5�O����������b��Z���wV�����H���;��d[0�i����Y���o�hѩ���/��`L��n���)�a'}@�2�U׌��'�Hc{�Q��R������������_�}S�j���� ���ekW�v^��'�P�*�z��M��~��$��f�*f�d[��˼�قK����E��8����`
� "�|_l�
@��y��}��9'��-YWT?�nh�r4��L*�}�N(k�%��#\�6U�UO�U�t�D�=����'�^��B��N��)3�z�����j��J&����Hmj��A���y��y�N�z�@������H%r�y-:X�-��9R�	q�U���w7|{	�[�"e������5�t��5"�/��Ʉ���K(A{���1M_�o���#F3@!Yp�t�NBO`Bo���vA���ɏ���;�����G@-��)�{(m,�1�3@t5�wq���O������V���B�R��,�#����d��֐0��h�>Y�(>ꔑ��KY��?��ғ�-v��R��W�x�?ń����;�8*ʙ��~��v@�-Iwm�,��9Ce[	�a��a>��=�_B�p��Q�\"�����<�@�|�y�Q!�gJ�Be������}�AZ �3"�� <��V1Q.��R�ށ���]m��X�k]�����:p� ����$��>�'zY-�\{�Cd>�b���jn�@���G2��|���s�fw�+����{�qD�Y�aбc0��k�es�����݆ E�y����>��8�S_�x���,D|�x`S�B�`������Zn���87�Bw<V����/=0��G��1%a���9���ͷ��H{RK��W9\X$�B%�)//Ed�m�j��YE��I�����(~�[&�m�$QGj�����`Qh��U_0z޼�u�@��`?��Y?(6� 9�mu�2�d3��ZK0>���5�<�iQ����yz}#y
pa�t���{�E%�7 L�]�GVv�*����R����c���#$��[t=q?��]^g��f���	����1��.N[�4Μg�^א�R��*���a��Y峾ʃ��Oh�ԥ��Z ��q� ��_Ңdc�1b��?:I5:��\}�ƹ;�'�0'J�q�ɪ��	M�K_��O#�2;��D�˭Ju��-�� U���q�=>�^�G1s֠��o�<+ދ9$��ZǞ^<"���5l���|[[�fi4fWU�:�)�võ0xw
��T<6Y�E\�(���H=̟��Ӭr�i�=E{<�Ԉ�/�#���O�������tTW'��E�ʻr�� �(MF�%�>��h���d��~�!�!�#[>\I�?������tؘX�r��Nw_.~��⤍�-"\(�s%��s ����j/>!���ȇcC����)J�,�k@��*�5>-��4�Y2���!�����ޯr��!�W2;|�j��e7�Hy^�ݖ���Ԛz�8ː�hH8]����[��x[| ,ii��?\r�L��H���c�vf�͈UWyo�C���D�;�^Y���g������f�:,kI9���Iѕ�@B\�wK������&lc�-E'C�}��a�o:��H��R5l~ѓ��F�N���%�0�b�o3����Q���֏ߧF̣������TYQ����2���03��y��:����"t��vͷ\���l_L��z����t���.{�'N�v�P�K*ud��r�;@4�{#X;&\/�Q����LΑ�;��"�B�	.Y��T���o݅����Y���Ƚ^I�|���K��I�
��$�̉�t�h�EVׂr�8�Ta\��lHJ�$&���:������is��͒���㜅�ڔ�''�kf
�b�(�'��b�*�.5\�h������{�ˌ��+-9�-��	���-?iͥ�6���r���F%��`�_�%J�A5�jt?��0�|�&�A^����JaT�����s��_3��DwD��M��jU��� ���1�d-��DP�U����A�9�?��yp��������і��2��59{�rÕƿs�'��4��q�@վ"j���!����l�wSr�6�iB���j�Ε�&N;}�����i�q����Y��x��wf�d.B'��	��P�n�zJ������ӛ�q_���&q����3��L1)�#N�"�'�6C�\�7�m�1=f�tW��l�5�|h�[F�Ѱ���������1�$�����Pg��l�#>1HF�#��'����7�`[��&PX��p�t��À�`���[0�J�/�25����A��Z