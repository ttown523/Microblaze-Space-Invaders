XlxV64EB    fa00    2c40P]m��
¿�O1w��T
����u�ڹ��<�Fu�B��+��(�=�������}�g���Vҥ�I��x0�P!qħ�7n�B�S�_ֱR�LbgL��C~��t"na^���O�{���Ԭ�_��L�d�"̝����ΉAD9�~pD?@�	F�U��f|Ȫ��:`���7��s٢�&�?#r$���}��~�Tߕi���`��b �=p��Ѝ�{`u@J�b��5�(�k ����֚��H��0(������ʊd�mo݇ؔ���33�R�3�Ϻ�nC3s�5!�q��]2J��~0�>ܱV�,�G'�_���+i�U(6Om�b�HB��c��W�7-�9+c����i��R�k�7ˉz�Y�ŢAf_��Y3��o"��)ŏ<~sf^l��NݑOkp�+�0��>�3c
�SC/����~�GԬ
��������z�eB�,�F��%�)�kڤ��nQjM&�a�q;v7;.��b|�W�b�3�xX��]_ى-��R��k�X+旭_�2�d���ҵ\�ϭ`o	��Dy��o� �n��1LȖ�ʈ�^�n���^d��j[�*��#��A@&�3(��`��茽?Y�Ļp��K��_ڮ�(�j�p��k )�֮���A�uo���ږ��;���&���n{C��H���6u�2v��Z���
�� vu�"ԬX����J#�
��b��G�	�r�5��z��&����>�ہG/&�`��j[�\����s�9��"��[� ����`�;d��C
v�!�e�&�;~\[6q���y�=�$�����Q->_���M����1��q�N����3��"x;(��qdY��@D�nV��~�/��.G�7:1������5gl��=�.'ϝ�mU@�]L��Վ;S�ݿ��vȑ<_��{���
��C�-W�2, �B"��j����O;�{��r���,��s�L��o�@}l貑�4z��@�2Ϩ=�=!��u�0�e0�r}���Yd?=7���Rj��΂��b���*��v��b��CI����9�u]8�j�dI&�S�x9;�%�5��ؾ�=��t�:ȷ[����S���l������Њ����6���ˁ�����z���#�GG��h� >���:}�ֺ+�+N���,�1"UM�<4Z�p�/��8�c�?P��<��L��%F�ta���@��.ǣЅ���Yi��g�S?�C��H$|P�g��s�N9�l�Y��V��l�=�έځ!��GE� �1��.\nu؉�au�'�Z�����Z�A^���Y^��ɔZ6Jz����A��l���<�ӖZܢ%@��Q�c�O���Ѡ3D'�Ah�oXw-�	��ʰ$h��nm���_\4(�l����'&I�^,�3��G�11�N@�&�9p�S&*팔��G>O�eЎhrV�Ũ^�VȻ;�?W�
vE Ŕrz���� ����5�K��b$�%}p[cW(�R&+$��v�S����n\��_s�_�N׀픻{�c'�x�=�o���wz�V-�l����D�B5�p@��.�l[D5�/��&�z٤� m���I7)���� �9H��R�j-�~k�5�b?X-[Ŏ���N"��f	�U���,�/�$E�F��h�5'��9k	��,�X!�W���!>
w27~K8���&�;���1����{V�sߥ��4�5�����A	i���7e��|��]K�!�
�.�a���@zi�`����\�F$�iχh.�������r"k?M?��}|0N݈��1�&f±�U�e��b1l��Me �`���u&�+?x��kuV�#7,ގ~�iI�	�4�D��v���ܧ1�����4��چ
 -ޑ ��Y�'�r�ҏ��) �Sq'�8#T�eλ$VQ{��M>3>�R��p��-����x���-tâ�F���P �)�MVjۃ=���P����b0�o��P�3<�VZ~��Y��%�F$��匍u�� Q>��1(��R�32����r�P8d �9�����|�ډ����p0CP)t�$��m����8���l�oa�h�%y���,Z)�o�ɬ:��� o�E���ZCu���-���3�a��0X�z���dc��O�d����Dq��	�x,�0�y��gf�(���"���lvF9cϤ)bSr�^;$@�Yq<<��'�L�<'���S�]"���6k�V�T�!^���z��
���nw-�^��1����Y����+qM�|���eW��'M�<����I�M��&�g!?[[������>�tuMSA_X�./j+)��b6۴2���H3����A��[ߔ�X�����B�G�>����];Œ9b�ϟ �WD!�e�q�F��
�1�L_�sp��i#�˿��G�&.a�8�{�%F�I�����a�d���')��Ξ��`s�}�A*�1A��^~�~!��<T��S�E-�� �f�'�����Κ橯�*>��;e!��ؠu�?���b��*����RPɉ�^�ݕ
[��������*mƒ�����ڧ	�P	�l~,n"T�:���e��ɦF}[�z�d��Sę�s��e�+�b����Ei7s�>~�͗y�I�j���l�t�E�搿�����<��F�M�#Gp<?/�/\r������9�}��_
݀JΥ�o�?<85�s����k��p�E�@7�w6.����:���	S�H�ų�k����}<v�C.
�+�BrHnq2��HXktk���*���0�Nz���d{�(z
$���۳f	H��<����G,!�eH��+X�0�0���q֨,��.��{�E�.Ok^*ʞ@����!��`�[֑ ��ʐ='�)r5[���wE����@��M(�(�ǜ�.�w�i4��1���U�������e��6#�"s�i�Ĺ�t$�=�ߕ�o�m�S-8�V���N�8<]���[9��&��;A��5%��R�a;c:<Q����+����ߚ7x�Q��,A`�TK�A�L�6�������� ��?Z#�a!��5H9��½�kK�q@�Jj���J�dnT�6\FO�\0Eu��
ղ�����JK�z�6q�X�U�B�H�{�P���"��VΡ}�塍�QC���f�䬤�����X�
�B=0TU�)���ƾ�TM�V�.F����j�}r�J.i��ܶf;�o��"9��		1?�KfS�#*���ʱڷB��I��ޱX�)@,]�J]AU�2���~��.� f�<���=Qd�t=����>�Q0h N��Z��i�ȫ ����|ޓ�������ݺ�j�����_������_"�z�6M�+��ܘ�97Ƙ~�B�d����.�y����a�!��rE�'r���ƎR7������꟫�I"S~����Q��{��Iq��q��Yx1�z| tL���g��#���4�{��6|46�dk.k�m���%��B�i_&�̙T� ��0D�m�IV���椴�
*j7Y����&��+PV����h�2��$�%O��p�C����J{��ueLsے	��Q���L��P��N�Η��6�"�wů	Ϸ�إ�o�����dV�[��Fr��x�;"h�Y)fAݯ�h��О�p>���ú�V�h"d�ߢL���YUf0�B-�v��#�9����a۞�n���ۄ��:'r8��{��1�N��/W��Ϯ.ܶ�5z'�yť(�ǁ�E-��:z۷��kޙ��K/_�Qor@$d.���ϙD�4s��l����&��@�6�Vϣf�[�=(��3qw��=ϯӿ�i�U�^B�B��`�P@�7)_ZH�aG��o&R~y����!���l"�HH�A!��(����{�a@��.K^Ŝ8�N~ߚF���ra�WH�8��t^ �i�v>�t��"'��F�̊��L���ӷ�6ͭh�.�w����n���y7�r	�r�n?��ѷ�ݏ�*Bֹ�y���6��Ο�u�ə�&U+,��?\��;Ǣ+n<9[�p�ԧ��/�D<f�I%|PŬ����u#E�>hІ`���vQ�:5R��=R��kc9ǭ�dm�X����gs��Y��C�����a�
c39i�l��UC��$�D����tTi�!�FzQ���s�ѫwӋ�r_�[ʡT8�QJϚ�i�}��fr�����q1e�C��Я�_�}�,�����B�xJ�q��_��0|ڵԬ�Ԓg�e��CZ)<�ʬ�ެU>�K3��VF�ٓ��Դ� &�5{�5)�ٖ����>?RWy�p�}����#�Q9ϛ�4�j�❠���(!��Duh6(8�.����$������nؐ3A�$��4�)���)�S��1fp�4-y^$�#?�.�>�Un����MxD<�.���P�+�����.�_�AsT:��v�|z%>CmVm�S4��bk2��q�/�(Ѥ�c��	���Z�Z��X���^�H��B�w&j���Lq��2ls�X|=��ل���\:9�c�5	��Y�C���������$�^��y��e�-��T$�Qȡn���:�k_[�Zf�k�d+���y�c,g ��i�b��v��s�5o�X���$�����u=�kƽ����p��pL�} �G��{��^�/�����&&Ţf����R����Ui<�B7s:+8i<y�y�wt�}MĀ�ѿ,X����4a�{�G��,@dw�#�.Pg �И��_ګ�J��(�L�����t�t���p�x�-"y�"4b��O�<1#eq��	A���k��)u���J:�Ʈ����uuhx7�ہ;Q�V����3�h�IΤv�f*��W_��?���=KZ�G�*�
F���BQ!F����a��Q�M�ط��}mK����F�T�f���+���Q��]�]}d�}�o�EQ�4�W<�9��ų�Y��E1��a�ɹ�j�Y������^�ՍAXd�GF �b���`���N��3we~�+6��W���D������	�|b6�/��./5���K-�gO}�
��D�17�e��kV��9]k�����e��@�Q��_��pY��l=�M��mpn'�O�s�0�|'�!��N�B8��t�{�V�ݕ��m(�\�C�D�����9�+�%��{kp�����-}�9_C�J�s�n�w�<�_�-\���������N�&��2$�Kr���C�{�H2��۶Yʡ^�	��W�������d{Bٍ�?��}dٜ�CT:�JCQ{��WiU{����#T��Q��σ��E34��%�Y�������`�6Ņ3���;��$z���,_�#�&dwC�jCaǐhK�q$֏�O7�>Ks���ʻ��]��I�%���b[-oϮx�c-<w���h��8Z�h�Y���-Lj�~��P{��� ��o��=��
ފ<���@C�y^ԭ�nͧϜ>6����n���0%���E$1m�đ��۔���.c���x�9$�����a���r0%��;��y�p�ۓ�T?��Zo�cl�6|�4@l�D�'�x��*A!��R�)�(�����U�X�q(��;�1��sb�?�JS9�'R�Qt�R��f$Q<Ô�Ɵ�ë��au	�1/>�1��j�J��&�JSS�@~@ ����f�d�5����=k�]�<��li�o�=.�=D�}h�*	F��%ϥ�g��%��Y��X��}�߂FE��Mf��F�<���#�!\�8�j���y1��%�:a�_�Y&�Ud�}���R��n�[6HJ�3ɒ�rC�D�Ń
��}`�8��sDf��F-T'Iz	Z.���%�a�|#�xjrE�� �N�r\��g�4M�+q��i�ry,��	�7�eE�����m��N�
������K�J�a%ԔW����>�hVH
�K�<2��ƂwZ�}�m	qf�q�+#&��]}���'ߨA��������<BNsΑ�X��q��xBΟ{���zP��dAx���1l�K�0�l:I�O��@T%@��@�մ]��ЀW������B�{��E���KA�����:��8O+�\.�7�񶗜w����X�l�)GZ�tm��5�����P�2��c��;�c�p�]:�i2oH�a��en���K�䅴�%Nj۸z���L��i'�׿ٰDNg���gkÑ�5 x~�̨p&�Z,|�b��k�O���@��k�����r�m�7r�h$`I@tH#���)E��{}Eyb�7�_�G���"�t3�%4������9��Z��'����TPk�]�ЏV?G������N"74sz��R]8CH��Z;�jk����{"��W���M�/e޺�.�|��UEC��*<Ϭ�}Y�zٚ�Y}P��U�*�'Z�� �ADFy��[	5X~v�f*��0��SZk�B6��#����J~ �1n��w>Ո��1`���o4_1̛ʎ���쏦��^��ɟB�:�8��)~�>�PV?�����v=�@k��?½,�P@1,ل���r#������`�����)zQ/�vMk���'�*��h\��ڿb`���cܱ����Kт���@�s�2P��LlS���d"��t��B5�%���4pV���AxV{m+�fs�����
2�}��;�J�ML�DS���Z���M���bA�~�Qę��ILd��M��g���1�D�tiV�k!�j���V� ��/W�碕ђt�mþ/��$;~1/��81�Xi0�K�FcJ��Cj�ő)�%����������f�/��^���n�p۳�<��}+��{��C�W�b&-�s��|�g�w��P��Lӹ\.%v��U��:���>�t�QF[?���@��i,��VV�ۍ�f��>0��[E@q��L�-G(���Q�U�ޤ�l�=���JkEK�Oz��?�Ud?��ur.F�:�(���;	؋E�*&h�E������JɔA��r�:?y�(g�c:0�z�^@+����W.���=�e��C#G���n��{ܺH����j<������7?R�@<�RZ?��5i�Pg�C}�vDW�<[��[���uGaoo%"5l��?��R�n/L6��:��~�b�`W6���:όó�h�P�~�	޺�+�����1"�I}�yI�
І�y1��N(��kO��3_e���J/zY�i�yפAS-;�u���A`�������D�9���z�cŗJ�bVu(��3>�j@�"���? �?��Ž��o��w^�nI��ť@��V`�勽c�[�����[���HJ�ӫZ'��@
Y���1Oec��xq&6#�-4���p���s��%�� �!��=���`���Zf�⼖�)Dg��l�N\ie�;��.��Z�kݠ�)�6D*aX�`O*p1����c(���K$]���$DM��Kw� �|��6	68�&ZFv��l�>ԥ�,����,���y[�债PvчC� 8LJ����V�6�O�{Xjm�mT<X� ���4�		{~<a3���wic}�j|h�̦��!�<Y���5yfr����o����q���G%�%������daKRܯ��T(r}����0U��E��p�\׵n9QQ���G��������3��b�T^_��|�6+�"�� M�2L��*��O�
˓��S���N����(�gzʹ�}����Jtɠ�u�R�@E��&/kW�I�u"R�(�:��'���+�䃼<�PA?����*�zq:�Rһ�vt�᫘�κ��[��I�J�%�K�q�/H����D@q�|B�H�P�]��<1X�:�2)Ms�\�$�v���y����1�c������u���Ӛ�(�\�S�p���VK��kk�g�b*�n�!���e�g��mW����wEv0�iE�q��4�n�X{�/��|�*��Ӳ��t�oM��f+z���4�3�F�����P�X$���@����4X%B8����D4��TKMO�͗ؿqQ�N��Z^�`
M�Y�k���7�9BԽ����..}��?A0���f��Ydc�3�]������M~H���dW�'�@�������v�0��:����_{���yH�d�n��,�>EN�.��q	~u)�]�wq%����?j���'=�4ι��h�B����i��>����cv�ɒ�7����5�q��7YZQ�n�IY%@Il�'�\��� �9���X��k�ZCvt���I���e����Z<i�(�.i2��B�?F�3ra�Ë>��U�%{{]�/��ĩea!�m?�#X����7L����A�WȲ?�r8 J2�h�*�Q�+4ep~z�w�VS�Y�I������6�M>��[7 �Y1#�t��F<A�ϲ!=�����0��m?��/��n����*<�j疿�%� ��v� ��/����?��o4�ҜA}FQh3O;?Ω�푩���c/��cy���FԠFV�Q�:������H��|9N�荪s�=/:z�$0߻��n��t���\K�)�}O��rk��k\���������N,v�?Z�$w	���G�|���=�G�@Hc�
�Mt�d1�՛�R"��kW��v����|5v�ǯa'��Wl�Օ%��G��7Yw��o�[k���՛����{�nP.o�n ���nK�bIYΑ��P"k���j����9D9Hg����u�d�˼p�:YײQ���'h��5C���MAGK��h�1a�kep/���V�=���z@v���n.��P��9�n{DzJ �R��O��q��l.&�j�@9$0�,j������YfH(�`*���׉�A�N8�`�@�)�^wJ��o���l��˘S�D�B�ɵA����߮��㤝���ڜߋ��|68�03o�87�a�ݓ��S�16d"CWԋ�׀p���qi�]�T�A�Їw��y[.P�������3@}mB���8�<�N����T����o35���EN4�J՗7��dt��6IU����V�gbΜ+��M��N�ϫ��UW�k9���dRY�Ú�XM㼷��P�\	�B�:p�A|�7�o�%�ɑ�}V�fn���מ��nMP��,;Mc�,�0o��<F��۝U�y���L=�1��͡7��1���#Jy��
��t�]����P	3(��EUK�����?~��+���_�I�/���?_+��N�n굳n_0�
B��fW��+W���q��/�<@�(89��F��	�GM�(�A�	K$8����]�����O�:��ZF�9���Q`�yN���s�:C�}D"}OA��T^�:��̫�AP�I;�QV��zܶp�Qh��z��tK�u�q�]�.YY�)�^a��*�\u4$���3���4y2�]�*B3{D������/yu�1����"��vPJ��&��Y0��{S؎�o~��8ݱ�>s�N	��Q�q�M34;I�9���_g�Ք����}.xϵ��n$\ A֘:f��]�䘃$c�Z�����a�g���2��
��9��j�]@���NyD���_Y�%u�'N���C����&����IUl=�ț$��T�W���F ������2ks�D�1�w��u�9$��mµ�7����/&}�/�C_{����n�����+��ɯ\����5��L�� ��G����_z�Q*q���\��Z�c���I�@|�6)�ү�HO��j"D��ёc�Ǐ���~{$����{�H��|�)�p��h��]�Ω�G�^V]�7
4�G,�D5|Sj\KlJ�������<�b�	�w4��j e�)x�.W��)��Qp�=X:��"�?�#R\�d����?g���E<spƗ뷮��ư��i�X�2.6u�-�?ܾ��ޟ/K%m�K,p�>�Oдہ�4f�a�H��3�{�信��-��J���cK�[��|-6�/�xӸř�V��D�d˂r�V/�vN�8(I�4�;��-9m�Ԏۧ�Zޭѭ؞�Mp��YS�(>�ګ���m~�R�C����#G*J֧���@�u.��)����F��5�#6����5��>^��ʁ�] ��TV<�VA��Z�")�M���d�u��t[[;.L3�a]3b_r�4A3qE�\Bm�k�z�#P������M�s9���J]rq3�C�Jx��F��L^
0����mc��K�8uƹ��vV��7��w;�PL�@o3,�����F���I� qbK���)@c��3�?�$�,���`�[���Ptx����eK�ۇn�L��`���T�L��y�XvIk+��դ?��}F�e�9'H	啕�]�e�l8tx�'���C��
�%�r-�|���({o�ʆl>��T�F��>���?;��zJ��U���R�o�I��y��i�7),:����.F��=�!�6�n�"�u������=��k����QM>C�� �B͜�d�1c����R�\*�t2LV��뢝�z�����7���݆2/�U!>A�j\5XK��-��U_����>�A�mv�{��_ȻC�/-B���z_��r o#\�*ec��c�ULv&���:���N�����"��-����t~��~AP�K�S=�������p�P��o��_H�?�Y�--�oĪ׋e*������Ll���W�|�/�Z�d^g���9S@}�H�J��1���-���:��lCzeML�]B�pl�f�_z_̨�`�����ʅ�� �!E&Du��t��R9����Fܺ�ycGJ�:�=6�?��\A �@k�̩
!k6���.PN%�sW'}�u���p�i{�9�.�zwD�^���>�h�݇P@�n�p	�C/�q���d&�9K�m����b�O�&��.m���n��Esl:�u�;�ջ���)���C�Q�ʏ�EnX�#VE$�5ɥO���s���9Q�����$L'�za�U��d�#;��jD�$�Nw^`<�J^�_#�H��W'eČ����~m�1+)y����{�O�?ޓ8oe!K�,�'�����U�2\\>L02��#��?�7r�I�hȈZ�u��Fa�y
���A����q����s�<�&�G��ݞ2�����E��l�E�<�J���_�r%U�6ۭ�>N��A�gueUxe�7i�!������)�5[-~Q��X�*k�'r�l��{r~����t�"�XlxV64EB    1171     490S5�=�*Ɵ������36�8W���ŠU���p�(�JC�M\Ő_7^�*�Dpsذ�K'$������0$�$B��E��ƹ\��}v��x��;�Z(�O����h�g"��*\���b	n�)�v;�Mk�'b�V�D�@�a�8^+��)�%\k4J�:���
�9�:�Q��aW ��]qMآ�g��u!ڼA.`P�+���K���[L���c4�n�׻ݺ����#�MO��/U�f�r�0�q7�kf!�]��O���2���6(��	m��mO ^�.�봆*���힭�~�W[@R��{�����4����A�ų��k�|��njC��\P�8�����)lw�4�!�F���6%�1�J�E�إn�\K��s|GǨEU���,�edWnن�JH���3Vj�x͘�d�p�3BM�8E�������F�}���d{������7�+�Ň�����Sgv�R?yi��W�_��$�?��уa�ǡ�#�놸�r�$%�����(�#���X�S�f�3�Ğ���>:H|�<IЏ��yOW����3f�Y�ھ���Q)TmP�M'MJ���V6�C_�O�f��������$����Y���ȷ�;��|� ��+�TwV��DA�.�	��3-X���3�����q́l^���yy�"/���!�L�Jl�J��A�C<<��j&p]�-�:�8�\���W�7MP�	כX�k|�l�28w���Y����m����u���i:�͑�Ҏ�$Ѻ�҅I!e������{�D�Q8�&���)��.�g�]�)kFL��J��b��bO�H�d�
U ]���*��~]������_}��m�Bx�TW�;q2���B%�_!�6h��E&󶌁A�z��Y&��"�����r��4��'� ,��r��uT�A�8\V�D�?��i���β��X��!8o�~�����N�$�y�AQ
�dc�ZD�[�`�+u�Y|� ��^y͟OC�Lw�ty����h�b6'�j��k�zUˀ|����O#�h�d���5ww,9Η�V%2s��E�VR�l��\�M����|K����4x�ص	����n��=m=�����'h�ܹ��f���j���q������K!+�lEhu4��"���ܘ��������<%�q���@y��$�