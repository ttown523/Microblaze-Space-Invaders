XlxV64EB    2e21     d30p�@�{�+Ng,\����#E�뢆��?i3��4R}R�J��5��Z�6
���M�Lˉ���*i�n���H���� h/I$k����-�pF�.��Ƴ��5�B��8�=0��m`�ؽA�&L�-3Mv޳�����F����Я��ͅ�E"9Z�R�zy<��s�41Ⱦ5*$k^��S�3�=W��yzIX�X��[��Gw(�4W'؁d��V�#�Y�NԱ'�ܷ����FDC���%����%e���P2��
�lS��-�y��ݍ�&�!�(^M��C�fAoM�A�e�5�i�(�n����Eg�����F�!����Rc�Q7,�B~�2�:0���O�2����h�JX�Dm}쉲�0z�V�y�Y���XC��]_���c��gk��;²���qqj|��ފ�� Ɯ��t*^�J��́E���r���m�Sv���,�E"k-�b��w^���l��j�M��l%���6���<>�pwK��s���8������{7�[��I
Z�����Z��\�Ӵ���+Qꐙ�9�'�@Lú���-�{&�M����#p��O�C4�ڃ>��:H�e���6P��.ff A#�a���s�#<��1);iՙ��o�9|H)Z`K����j�����.o����!^_o]�
0q�T�I�"_YNʒ�����s�]��Xآ��Ջwm��%�%�g�NDx�;@=������"0m>�i[��_��ɲ2��T��ס�����U�Co��x�I[Ɉ`�U�p�7�`�>Ir�N�e��ra���a7m��;M�&PO�V�6�O5h�oPa@�<�x6�LQ�^	�E�)+�s�z11*�@�B�,��"(
�+�W���J�lg���0�.yMI�q�	����J?��.����EU��/g�&�n<��B
'Tދ�"���Β���r+q�RVhO7�>[E�a�X2v�>���bE�蛫��(��%�D����IR�b�^�)�TU�����h#��Y8}k<��� �)Ȋ�;[����옄�#�8U=���������bt'�0G�wP�R���r�z���8\+��w�
�Rm�P���i�ywi=A�t'��x	�7\��!�<���*��]q�Z`��Bo�ƃ-?J��a	�n�]I8�I{�8��'�ޓ���,�Tskw�$� �K��� 9���ĳ����RD�O��S�|���D|�'��_m�!~��yҴ��j�]���d�;'��������)f/��i����St� �ɦj�re0�$�qJ��8i�h��L.��Ĺ�n+��j~C_�������N��"J�s�u��� �E��f&9�ۘ)�z0�ף4l�8���|Nz܉]_Vx��$�r?��K��_t�Z�R�j���<�,�|=�M1��=�;��K��l���ʨ2�]W(�iDa�D� d��}����']lg	�ꨲ(�`#i���$�����u��7I�7� ;넋udl���ړ�a׶t������,���y)�<�����������d(���MF�����UlqA]k{ω=k���2ν�.�b�>Q�L���s��9�]����8ď��ႊqx�s�����B�j�˲u�|�w�m�JeN���<E!Ր 㠕s��?�X�\�4l}ڏ4t�굳��Xn�t�/��RF!����[�D���iܥ|�D��ݨ��4�`�k��>��1-�Ѵn^5�;H:�HY8��b�[C}kLB�=:�SIk3��^�*'v؇�o$V9�:`�mH��<�6��A���L0H���R����Gȥl
\���cK�ZRa����
e��Ýٕ!�T�%8��n���\*��#^G�b��Yq�܇3k_�N�kb������N���sf �ph��ʐWao�[�3Յ�ظ��'�w8I�H��������GIbw϶L{�q�U�TI"i���2�ܸ�}Z�J�����B���OS݅[��M���4���\���7�8���B�fF�������J������Rb��͝��ݠ�!��y��z�"�#0�4�Lp،<�XI\����#��d�aaj��U����a�Ȇ��g�'����ps�թR�eK������?����B��&�x�(P�hO�de�Oڍ�;��Y�C�I�z���W��D�bjV��K���/L�#0�}���BR�ul�gB�r������a�W`�
¡m%�TW����m6�8�P �N7�}�J9��/�%.�+�xR���?�0�����r��A��@�Ƒ���?Q	�!d릍���xs������|�����t��0�2ɑ�/ c<F�rŉ,�Ѡjۛ@-��:���Oɔ�J��ġ�H�È��0m�<�o�C8n�;gR:�#I�>V���'���t�J<�^��]_���ȓ6�Sz�Ӆ���#Hz�6���B�?�����7*�>n3G� �n(�I�9�USy�?���jw�{`+���=�p;����l	�>4������O�s��'��㊉> %/����MtF���i]����W�:��"��̺e�RG@R�!|���`(o��_c��뵨��e�/ϏV�hB ��2���ZGt�J�qP�!�lSS;[ɦh{o=�ܱ�� �I#0��Aͮ荞B
��p�0�Ж\��\gv��oH�-7V-�ޘFMY�;�J�c�k՛*���*��I�kz6>7eS�d�ؤc��on3Q�S*dr�����pϊ���!�%f׳/Ȱ�� ���c�.�ۀ�^�@W���ϐ4$E���i�C~�y�U��Qͬ�L'9��ˁ�s��c���@������`{��Ւ���G�c�y�;����Z�9�/o>s�Ӷj���O�]��s��~�lw�˸m㤰N��5J-n��|�S)���Qm7�,F��k|σ���t碕��iӶ��ũ�Id�)�x��h����ɟ�Qj�������U�F�-�@P����=a&��a��hݬ������v�c���	�����t�:7�L��rw$B5B�q�j�R^P�1&�kʓI��_q���-���=�cb8����F\(����쯪�Z�Z6��YPXMbI%�����c��4$��ܟ�X�P�>��0�}���ؘ��!�+��vt?�V��8d~��g��;��;G�K����ܠ��eP���u��j��	,�<ad�����+$i2so�h'���ь ���� ��Ͻ���!);m�b�7�ә���`����,��/aG����^�	�|�%��[�r�h�*#�>�?�����-�0�Y5�Z�,�
f'G�߱�$힠F��� �;�H޾`j�9�!