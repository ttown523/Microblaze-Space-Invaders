XlxV64EB    a7be    1be0NU���?�"�S	�	S@�r��D��q۳��:��e'��=���;�y^L��&9<��}�BHE|��^���wm4�{���x����Ra8����n�2��]/���!%��0�>`2��1_5�Biр1;u7i�#i�~¾��(t26+	�Wp�@T�3��J�v'օR����BYxP�Ϸ�&s]f��H����]����],W����5��|;��M�? Y$�#X���u��n,�2nS�4pn!��!F��K��(�~ʑ+0Ѻ48�a��y%���!���g(¢�pL�x�#cn<��պ���ŧ�������u��.|�d;K{�{S;��s�Zh��s�|}dC0����r��'j�Z���݉�9��$�m L���+t~��Y���6ܹ�{�$�;���R�����eU6�w���q�].n���%�3_�G����w51��.l��4��$p��r��_�C�����K�J^��r���K�tnQ�o�[����tl4/]P��a�;X��<.gp��Rj��G�}72�s�O\>�����V��S6=sJ��	^Q���ɬj���s*���5�v8�CP�KB�|��/Y�SDqCYE������q�W5�z�H���`l�^����X�`�U������,%ȥ}�*�r�Ϳ_�H���JwP��0�������)�zܣ��0C�j��z�K��^�ے�^'\�(�Q�/��=VnG( H�f�V��o)o��Z���i�X��H��T��ݿ��?���;CVu,q�%&!�5��x���O�;�ߊL��U���M�Xӹ`�(ԯA����5��"%�:�h��3S�������W]��ð���Oh�咏�2@�Oo́A�Å!H�Į��i���PFߵ]hw(�R�]�B��(�ϵ�~(y���{?m$�%�AL=�[��T�t%!�+Ҝ<�}CkJ1q�t܆j��Lk��dYB�$A� �-��S�~��M_2	VbK�ErG~�����@�_� �<pU��kN�C�o��#�w�������l�܉_LJ�kY�xᾑ�A����xa����M0�G^�-"���aR��OVT_��I���n=+�R=�2$�q@�Z�a
��S�tU�E�r��d�U�V�P�f~�"2H��UU��� xw�?{�SͧAO�k}�����ۻ�G��K�PV�Z�c��,��Ĥ��Y������`��*�'��rt�n�����u���:�oƽb϶�$�@ޒ�Z�L�6J9j�k�Ծ�dƻ�ZQ	��q�kz��M�I���p)~���9�9@�c7n��[/krS쉀En:�CG�qȜ��W>,p��;�.p��M�6V���{��[(���poX���"�(�V���$��r�B4���D�(ڟ��n�\�	�%����/U�����S�w'"��X �����rò (� ����S�XW'f����|ʈ��9��V�R3���2�	x�r<��B�4�,ܱ״��b1\ޏ�I����W�:3�5T�3A���@?�:fT��E�(��=���|�Kh:s�e�)AͽC��r?U��b��ڀ@���Ī7��svc\�\��S�)o�B�Hw"O����"�B�"�����0�O���w(��{�`�o�bk�@�>C�r�F��jc�q��wB��}Ih��׽/S��^�҃π�.�
�(h�GK�^p�H�p��u�K��f��c�Hkq��+�\�%kv���4^G!�5�ڛ�e�I�*�R�!I|I�B�f��$�S��dRA"`��,�d8���<&�h�&�C���6�-N��)f�,�o�x�N�f�����X5�JB]��� PL�6�Q�-c�A[�!�#��+9��钔6��E/�˄��k��:�A��x;��;�+H�+jS-m��2��'	�\y3�⥫��sj� �B	�v�F��r[����,@Wo���i�{��bQq��Q������C���pX�����HS��u����Ĥi�t]�v��F�U�혌=xd��l���3��<+y}31H�C�֏��`�Y�DK��ɣl�6��@%�V�b<N(i�jֆ��ᕫ��(V�sϞ%]C����[�3����#Nx�&��;k���\�*��'��ҷ�:���<�6~�D���j��3���:9ᡜ��䌎:�vՄwT�V�G1�g��e��g�Ra�5uH[L
L�oQ=��UU�z$�np�U3��_�o����)VS������OT���w����xF-�T�N�c<�6�˰���p���8��m��G5@�!�v_�>�*5�з���e��hN)�t� ZIY����n#:"�NC�z&0��.Ь�+"'�D�
]�Ř��P��9q$/�ॄu�ԇ���zNY�:�{�*,�Q͉�5�	C|�w���>=��w���Ǟ�[���q��iL�-C�H|��:6'=�-���:�k�6wő��q��&���s��h���[�R]�ȂH���F8�*�P����X�xgԄ��Oi!O*KM�̔��>�M'�D��PB�T֝sI[�o��y��5A.f��N3>]}<��;�1��D��M�8�v��!)���<n3( <�]h���R?%fA�G�1h\��[��%e�'$�ߩ1o�q$��^�'����AL��Tiݙ�{�u�A��N�AA���s8ĒЭ�uRz�?Jr�r�{�R��̛"̞e���x噫ʓ�c����$�i�.����O�~��^pn@�D��:ɳ���]���T�a��<�s��a��߼�7�Z��u�K����5L���0%�5�_*N�喜�{UIOzk��Mh�CA�JΡ)C�J\s;7J�e�_#��S4����4+�;����}>Z|����,f�9+�S��ʟy���a+II�s\���C��5*���9�0��rhYհc\"��B��k~U%�y���{�R�?�v��5�܀���p�s��?TY�����,�+��10�� ,*{���*�f]��[��09E�m)<�^P#�����`(l�k�����vC螯j��;Wn����DX0�0(�,�|���/O�������i;����E���ôh�]h�Go��R0;8`iG�aP��z�`)��םX~�Pm�D=u���6�Yfڶ�����?�����*��Β�.~0��FR;r3��f��?�h����ݘ)���>O,M�伋eD�=�&TTK�h�m[�U������G��CFb�#�J��׹�(n&{�
����k�7X�c(�U`�e]��B�g1e9t"�1�l]Ǵ}H9�D:��=�!���T�&��S�Y�y\�ʆ�Egk%�����;�B!�ˎ��Zq(C44^	�"u��D�s��w�s^{4T���W��i����k���hZ2s1�O{���#��< ��?`����]����L�����.��6�^"�y��������k1���"�܊��S�@.y1���w|�B%���2t`�F}K����*�=�YK���+��
��nH/ep"�e�_i����������N�7a`���Y �2B����<�m �Fϴ@���A#,Hl��Q&��O�UJ��Le�̐�"/'��܂
JU\���:=�Ǝ�o ��{+��a���mNY�-:���~��]��I�_���_�ZW{:�֦��7�θ85<ӘH�'�$2�*]<�f(^�N_�ؘ���^���3z��C>>�� ix5˙�.?��U3U��5���w$�9W��ї�ۛ*ħ��ഞq��v�"�Sn��8�Ϳ�F�� ���Ȟ���B�͔�&`P�vd��:��*y�ۋbV2� ���(�F�1�N�H\㔬54/6��� \e�LWeKn/�P[���f��W�2�Pil4�� њ�uv������n��D��T$��ŵ5��	(=�ޝ�F�r��wm?����d,�AR-�����%��$s�@۪O�|ഋ�g��i�Egb^�BAa�)��L$���h~]^=��=�=j�����X�~%����+EP�1�t;�W��u��A�v'��d�N�$w�_��X,��"r��ۨ:/G 23��E`q�H�Nj���h�f 3��緆�	�̫yy�$Bld��>r�p��e�A����"E[�Q���_��&}-�S����n�Y��HhC���p�E=�^��.ِ�L,�H� ���-�9I���n��4�S��?/ʴ��08�{8������v:֘(��LZ���RҜd�U=>#.%'8U3��N-���t�cd2 <;�s\��=y�C�q��Ѝ�Y��@��|f�z�/0�]>%����� _��Tخ�c	
K^|�w�� �X���E��zߺ�ܩ���3Qԑ3xe}���+{hn��Y���4��gk;3�#�����]lb�P�q;��f���Z�xc��[��OB5�(��\��@��ڔ�ٖ�v�ɾT	V�[&X��%sA�z��W��B �/��ᶳ����X�7��	��r�X�sGD���s<��io��սm���
p*k2a��P�Ϳ�rٍ
��iL�����$6��kL�6�WO�q0ןG��/a� 7;}Wz)�W����<��Ù���F��kn�!Ь���^ձ���\�0^�eޝL3*�!�R6t�(X�!c�2:� ����wx� �_��@�M!'�6�n<���xV�������޿��][BYrU���0;KXIw\c����L�	�+c��ԙՏ���pq����'�m���1J]���^#�K�T�A9�QF2��9�u��*fо�z��ƽ�O��]L-]q)p�]��W��4c��Ǚ�'b3\[�B��|��|�!RA�u>�G׿���``]N�x�-�:9=e��F��!"s�Na3�ZH�W�0������|�uc���<g�4|���(�9{13�4��]M�J��*,���s�c���{Ak �wG2v���c��$���n|��tE�����	���5�l�Lwc�K.�(6�O�'ϮD�c���y� ��!���6�G����r`}���@�����L�a��i�	n�(:�Ѱ�g��#]��>�p��{oۘk�=�宎]��V�u�'�\> �2��\�~�g�7Z�"\����ěBc�Q�TE?�n�nc�,�yޘJ��Bm/�qI��V��/}��?<�fji�K1�L��9X�ǞSrV�M��G��:J��
Ƙ�U��4�����EES�������e��j�L�e'�U�R�{��s�n�Ƣ�p7���ⷼʺW�ň�[KNp�V�#:h����$J�W�:���(D0 ��)�A�[0��ؑ����(�<�ǵo����;���J7��Җ�LU`2�Gh�6�j8f&������
�#�vm���7�����c��wbOQk^9�")���^5`�ӏP�K�K��r[�sw)4˛�=PQ�#]���y#e��q����������q�t���jU���-�yH6R1��ܶeUí�Ϩ��=)d�=�^�,��Kh�����+�Y��a�Z�2�j ��k͍,��ksd8#��˹��ct�RM����gF����u��0�e�ı�D�_��6`���[!w)MtO����mЋTr�j:���q�T?��mo�'�يr���i�g�?�����ZJU	�o�M��OkV�O�Ng#�e��;3c���㰟�p�����q��n�i`��p�V�a����&��nb��#�Sv��3��&[�&�%�R��, +����dDA��]�z�:or��Q�-�QVif�a��j�]x\%�<nNМ.k�D�bq"�v��2�<��$��2S\���%�0��Y8�X��>F����h�	���ɒ�拥�?`��L�l�mu#���(}-ж�k,�ݨ��mp"�Lڡ��b;�Dc�8��h*F������lx�}��Z�;�]D �lY���p:��kq�l�.q����S��@@���� [�l���<��A�����u
�<���q�k	v�>0�ܨ9*sju(^���V3��4��|b֥i�5�.J�o%�+@O���
Xx��@z���(����Q�Y���s�]\k�����wr{u�Ѱ�ަ8I� .R�}��g�A�tw�=)ؤ� ��V\�3|�S=F�&R1��s�����Q�.6Y�#KQ9�V~c���Ί���F �4)TVU�����JtU���!/5`M��`�R���G�5j�� ��\裛w�#����V���]~�qg1TxR����e �͐]���$�F��~�^��5�_�VaK2��ķu0�!��!���
���ni�q�|�M�ƞ��M2yPO5��$�jxFP�RqI�{y�ꏈ�߿���\B��XB� ��ѽT��%K:^X3����>L\@����B�z���J3m����F��ѫ,�#�}p����5x̯ͅ���@��a��3pH�WTX�$�GɴpѺ��T_��.K�V�u��[�[���:N2�̚���/���ia�4��"���m�JkƐ�4���2&��6����]��\�(_v�Fx^��8�\>x��a�ؙ����H���h\�wP7��z�ct'K�E��kG�^��@=���O��} �v�:�o��N�D܌^�KǨ�?����G:[�3FU���vp�q::M.�Q$�'MQ\��0L$�uNx��摹S��f��P3���i���n�@{k��gAz�&�؜�'zE!"<6�HpS;���v8ܝըH� ��
R5Ռ��W�P3�6�O������V"4��E�)�"24VB���� h��� \��=��Y3R8Ei�>�]��ip���~�{Y�B�l ��D�zP���x���$X��rd�:{U�|�^��O����-���Ƨ�&�7�ُ���{%��+�d�3�D<����pF�| �(�{x*�T�kwd^	n��-V�c%�~�d<���&0QҢ.�^��g9c�x����xiխK�>y��,�`U�	ƛŇ��#'Yi�+��FŞ3ac9\3���lDM��