XlxV64EB    5648    12f0ѻB3��ҝ)ave~�K�5�$'��Sہ�{[��7v��n��sׇy
u�}Wz鐗Q7�������:bQ6��@M8v���\�:ơ�"�F�����C���<M܇�aRaY?�	���^vvi,Q��~�}��pLA2�I�;w����m�}���~4������a�qs�Tr��o'���6,��$����Kq�ꘋ����^�m(ʡx1؜���Ey��z�l�P�ۆ�b�>�?�S?�!"�dȤ]o]�^�N��_vp�����u��X,��PFJ�=�,��"N������ +ݯ[�H7:n� �<	|!@�+	�MB��9�Ҕ�1m��y�6N�<�e�̳����&u|P�΍"2J�v �߰��yQ ����}�_[I�N�!Y��|م�S{�S��gRr�ډ�Oi�\������F��Z���/i�N�1A2�W�;�HZM���z}��\��F��ޒT-o�]��Zs�J����{�4�R��C����EO�D��H�Y��c,X�ᇠV�ch閁ӂ0��уѝ�����D?8��Ɠ=\�a��I��Sr0/V��Mt��T+M+���[�pI�ĵ�$���,PU�m]���NÖ�Ϋؐ@"����o�M�!:��|\ٻ�HI��*`�dX�E��Q��򗴐����:�=ESe~]T�!���P��k�毿��?��z"���)ku�~(Fn�}s�5�1�&f�޳�4��˧3�l'�+=���Ͼ�8|6���u���8����%�/M����p��z+V�3֟�/I�}���#92�#cZ� �]��bO^B�Ivtx0�f�n�K��Q<:eՁYӅu� �9���D��Y�Dbɞ(L
�s��
�m ��n�0	7��[^��V���ż�!(02��N��o>mfķ���ɩ��d1j, K���_B�\������j >{��;c���O��R��@߄�֤�O��G�w-6����3���kPz9�	� ��^~U��PK��<��y���*x�.F"���f3S�׎Cx^����I�{0̥�Ē�Sړa�XjA�� �'K�T�̀Z���2�@'���oȿ�D\�-"��x҇6YO�Y8��n�m�`	^�-�.h�	m�J��=�U.0rI2��,�����#8����$����f]\W�>d�g�C�s�8I"��a/��G���F�1�ݙ`�،�1m�]�7�]���R@��퓫�f���O~N/b� ��n0ی�<�Ί���&�&Pշ����ca����S`����ҎŘ��FcF}d8�^?�G=�	����g�%SY���{4�{�-b��.�3����c���'�u_�~e�:FQ��6�u�F�q�I8�l�(	���Z#]�ݠ�*}_
C=I�gWDU}��\E��W BmIRɬ �O�av8h�toKA����]�>˾�1�s�Yl�0��"|Z(��@�P$@i���BJ���FZ�3�?g�]EpnQϛ5m�D6�]�N�rQ|9~إmy�G��|>0����y8�٫�+qJ��u����~�s�Cّ�pR�*ZYM���a���b. �$�Q�o�_��"�M���C,�3�n�V���/-���q|K�?�;�-�\E�T7�+������ѣ�tHP����j"�q�8��i��6T�>E�l�ۼ[�U�Cb!	"��������HQ�,j$ɮvSoED`�(1�S:<8{�ޮ�����X�)�n��¢��xY����h��������G���N(v��f�"\����J�+���P�=��,�=�����R�op� OK��vO]�QHd�E�ј�Y�A�'ϙ��X��Hs���E�6�At���1'��ۋ���R�����0�ɯTJ�� 8k��]�[�1�2���C��Ԫ,�AO�3߁������,�w�u�ù	�6p=\b���y�XdQ�4��4���fQ�bxYٱ=_�Ԫ*{|*7�I_�K���6�2����:��4��Z�<�m�v�_�9���Xl�<^���R�f�� �eC��F�� �_���sF���>�@�+�]�p�햢�k�\�|�<`H�T1�ypo�zj��SNV�@���oW���
s�
FdhXUY&��L�<S C�}#�E��s���̀�$�x-�F	�����A�Qj$(��:�y�Ӷ�>��Wx��B-�zq2A�GlX�B�W�� e����aߒ���yO��Q��=9�gƌ�ݜ�I;�O�<�1�F�ow����|�7��@cÏ�R�d���s?(g���M�v�.�\����})��)���!�JWk9rѱ���X&r�_L�;kf2p���	?J8v��8-�yڀ��t�fxx��)��]O;�.@��~;/��Au�7�[�2� u�\9i�!��r��C8ga{�^^����
(�a�i�N�6�=á|�v;la��T\�T����Nk	�2�7���F�H�#�W4����ǭ`��4�s�|��9��\O����=�s�[�-�Nt�<y�QW���p&jɩ],�!=]�3���� N����ق<�D(ȓ��䚊Z�/q�Б��x�Z�V~����gK�#��z��?�1%���.��%ewߊ�`�[-��JYQ�J0(r�˃ڸѱ/+�ɡ�^\ͭ���/���NJ��A�z�H��/�bI�S�H�ڴ�B�`|L$�bUU������{�J"���*�ۈe��b����"�A��3n����-� t��3"%�w����:_*����ᘡ�X?W�0��1��&ԞԎ��਽<�+�oAP<�{�D|$z
�_AҎ�섏� ~���7l�_�a��Q�͟�BD�c�d��*ٶKWK0�n��������5w|��d]|�U�i�0n?m件��V�D/B
�	$��`mj:v?��8�m.9��C�7kg��vY�&{��ܐ��<O�Tq 	YRg��":5/�A���g54σ�pB])��M��Ғ5���#>U��+��]��> ���RǷN�b�x�}�$���@� wq�P��{�@��5]�0�,�ՇP�R
���I�#��/x���-a���(�^��D�e���[� ,d�L�J�B�^5e���l����}G��<s�kڣ��d\/�,J�E�_�o\�э>��H��VFA����N E��o�:Τ��z��C��<��:��Y�K����l���f���F�Q���W�[��>�~9T�|4ʎ��/�O2���U��q�Ȫ�-�\��Hd;��A`���j�ٚ(���
o q)s�1c7	�/���6���@{#ߩ��6A$Y%<�~8��8ju�D��_9vY\g<iq0M_��0��`�xF�&��GH�/��y�:1�pe�����6�,Ur��1��"��H[;�8u�N�ŵШ���'r��E�1Q��!hV[_+F��ǲ�6`�9G��ۊq#��7W#&���H��wj�J'@�32o�h9[����PO!k�((vqඟBq�2��Z��d�ˆ��hJ{,=m�~�>=��3��s��\_���	�9,�o��S��AE�����Ť:L����`[o�y�Ix���4{w)����=;q�B)�p��'������(i���Ygt��<R�1�m�v������`�a��N+�	���ǽ<q�	�V�^Fq:�`e�Qf��M블��Rv>���0>'W��sE������ pW���]�W$���A{���-�1�%s���e��0o̩?�:��'ϘW%����z�=w!@�[y\��5� �3��u���\u�3��3�l�X=�T�g�d���7wq}��L=�A��?�~��r���[NWg��jK�Pۡ�ry�
��>�����DXu��I�4�4]�W\�u��Տ�7�AF3�Ĭu�F��}�T.)"޳�H��flj�:�9j�>"C�@����u�[�V���j�����Dm@��������!~Q6+ݏS6� t�8O>���u�9�4�ѐ�E�[��YP<��8y��l�}�%�e\��9��|��q�G�"�7�ef�)wh*�ڦ�xz1%+������F���Ɲ.�+3-��gv�ъL]��/��Mp��M'�m����22�^�_R�:����/{�$��c���|���2U��PX��y�ـ�мv~��c���t�!A ƣ�~* ���}�&�"���*0B��k�?���7��!���E�Pt(���
*?�(�&A��p��	�5���|P;8�����L�S�D[Ш��䪛�/�=��� V�w����J�T�2 $!_E���(m�+e�Q���%���Y�����R�D$�M�e�#�6�ہ16��L6�����'T�M����a�zO�K`zN,Ҡ�9*p��7�g�S�|cImA˂|���@���I�V�<�bQH��Z㺯�A*���"�/m������DŸ»>v&�qu�Cs�2�4��"v�]e��O��;[n�*Fvd�vAHQ�nDm��x삻Rw� ��ML}!��Q�~0���t�:�i CC��y 'k1R9@F���H��_s���]8���ٞR-�҉ʒ�����T�������bwPL�p�RA����;�W���b�, 7��UT�͉�3N���oͶ̻Yү��U�T~���R�k���C���5� :�5�������Ɛ%��ky�f����T��`��Q��}a�����s5�19�;�������g�
�߰6����{���?ӴWպ��M��T�Vv�
 �u���XYDZ�W�#�[?