XlxV64EB    2a48     c30ˍ�����֖XD�=�=��8z�۱�2(��"8�
�].K�^oښ����7��%�Eȑ<�qK��(�z�ȥ���Ap�7A�����d�_`ؤmЃ�0*�$�S�jq�W����{��pT�9z�5I�;��<ftě��_�a
�>j/�x�֟������b�������y�������<��ݵ��J�m9�1��-p�e��V{ �c�n(����>E4���۔:���"�n1�גö�K��<�����Z�������&��t���2��Aj�$pE�4��͈t�Y;��OЖR�9�{<�_���5�e�+{=�e6|�kO�3��M�2*
���˳4�[z�Z�ҷ�<u �O�����ɯ3�f�:�d�|�G֟G#�4�~���\.�cl'HJ�P�N��;L�z�r�U�`�a	�F���S+��o�:��Am�����ʿ����#M��BO|A��g��z�9�	;����Id��C���ިT�k����N��,^�L(��N�5՗�:QARP����LOSo�ɥ\]vKY��A�$y�{,�O�����������PZJs��U�s�_�v+�61�k��ek����ѧ�50}�F�I��c�!�Ń|������o\�Z�xGI~�}Djҕ[��ͫ�,:%���d[��/�M$ߺoH�W�X�c �/�4X��.KnLwʝ(>��6NicS�w8� ��l��� �j]�v�5�=��h󪮑K)�)si>:��烶���'�ƪ����?��.�D�'�xX��{$��ƸZ��G�#��A����7to�pp�8�d��x�70�b:nA��hbz��c#{�TzӲtG4_���l����Nq<ݘ+�џ0��?qjQ���0�����)5�� "�]��:���~��qU3�����A=�$R~���9��8����J����q����BH�h�IYc:i
��yE�
��MJ�^Q�u����K[v���qº}��RS�:N�����p���H�)�M�I<O�5o'��y��U �u"k���w"�D�����yc�+U�lc0<���:h+��ő����5Wj�0��:�B�,z���զ�J!��gڷ���@�^��̓���ln�R��E�����ti]W���e�Q�CSȳx�}9Rh:��e� �l3��Q�w(�Sy�g����ۍ5���B�H R�&.�t�ؗ�� �*�l3C�Mb��-������zDߝ�XD #"��1Z[�0ӓ\�nB4ϳh곐z5ȊcO�>�KN���e��T�,���&���I�!̅V�<��v+�u�+A�ֽ��45[ 
�E	1�_��aoV���r'�k��G<!�U���\H �۴Θ�S�m��L�����`����7ķ\A���d֡eB��ȼ��a�;BZ<a4�R�������wluԦ��y��i�(�߲)��&9Bg�)����*��aR=ā�����[j�	s���s%�17N[�N�L��՗v6�~@��έ$$�D�{:x�H��r�{�A��f��<l���r�]���s��/�i�Jf�������2���Cפ��d�%��@�,Y�q��@���61�?n����\�?���@�\�,:�mh/�]�,�u��NJ��P�yg��¬�8ȣ��2	&$���#4�'@s��r�[Ę�͇ѓ>f��[�[��&���@d~:[^��F�	Ց������X����%��� Y
篲�AA+
nl�H!.Y<;J1������ǡ�h	�(g�[�}����e�p<R��A��i#&�鼢f��v��X���JP��Na�X����\u�	�٪�?�20��؏2&��������L7��(�������=#�Zo҅B���|�ZD)�	��vo}���j�+^�}�Cd��{VͰ(_��ͷv0�<'����c��;����!!�8z����UB ƪA �.�~�PZg{�R����V�p�*luX�-��\A䶲�a��-0�%�
���sO��-~š$��㇊�DWiF!I{�[7���X�D]���.�ҩ"p	�̱4l�&�;�l��J5r>�ߍV�L孶��lP����0]i������4�M�����M����#�y��y�}�=�0&l�q�;�޲�t�uCUq1"�B����jͼ��L�1�QK�Fb����d&��Yf2c^C���,�74B�ђ��,&P-�r[Bv�)w>��:��dTל^7����z��ix�:e��^���:[������-��j�4�W�����(�nu��vf��C�����Q�{Zy�GH�@��kc���X�i�g٭An�H�"����T5/p��#�ՊS�2 M��|�ar�J�~j_b9��g��i�P���}
{̫W`Bo��z��,B���}t%C�S�5=�RHԳ��:&]��;j��V��}����g�t���B��_����5����T�@�?'n���1��6�u�Y����g��V�1�sT�>�Q�JƗ��yXT��XSJ����q���/��{rA
�Of`&	����Z������S����	������|@�>��͛X �N"{M�{�5�j����rP無�鋂���yV�p�u������'����k@̻�\捩)N `[/$ʞ�N2`�D����%����t:�����.#��"���+H	9!�����r��.=��Q$;���{�ή�����`�C�缨YNx�A��B��\�B^�.i|J �h�	�_/�K]%��~n��k���=���v��P�hS9��6�̬`@���Y�1R[cud{��=��B��L��|M�5|��ͨ�`�*�+���D6�N�*Is��h�je�l�K��;��z�l����φ��8.�c�#�o��P�r/��Y����FiE���w0[θ5'3�B5�,@tN�~��b�X)<=<�}%�L]&]"�����p��D�>LxN����)���R�x9��6�x�EcÎ�:6>_�r�UL���]������?����ņ��*�tㄭA\e�	NЕ��[%�M��.E�֣@f0��t�R�	��(2�,��