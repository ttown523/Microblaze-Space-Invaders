XlxV64EB    fa00    2e20	�*���To�Դ����G���b�i?���#���,�\d��~�w-�E��0:ąO��nrWh��p�5�EZ�+��ˢ��Νnu��Q]s v-3y�S�����vV<�nA�Vm<ZB�S�U�����q��Ld�Ɉ���oBC��@7�mנfCJ�X��k�<��"����b8�X�f�%bk�@7��66��W�E�ԁ�?8�����k��/> ����~U`�es[��=�ܿ��f".�-��}Nm����9C��<��NU���ԋ�j�A�S�2�qs�������7-��Ͽ܄��r��&�^t���y#�<R90^;w�i�p�U�JzJsP�꨹���,+����Y�,��=�#/�;X O�0EO�e묻��e3�'U1�Xb�H�͛��/�YM�ve}`������f�]�v9,�2�4��=C�,m�C���*�����J�������!���&�Ĉ�?0�p3ub�R{�D�0s O������^��־�T:�0h��:0$�0����h'�,D��W��\E������������J�i$"��-`U(ځ��%�C�e��*_��;
.���H�#���	<>X�����`=?Y��'Xpv"��#[X���7�Ԝ�3�'�c�QJ�Ԛ	��;!u�_k����)�Fv^*Sj�x�֟w����Y�O?�E�@p,qֵ{������?h�֘<�6�F��Ar�+��_��H+~yҵ�o��ů�?���J�U$�]g��ꨮa�C���k�;��m��T%�bU{��'�W�1J��s��F��
��F������4��-��h5��B�Ҷͅ�\�K��N�r%���@2�Χ׽�O[�rtI���V�C��x�j��>��p��9_�*�aI��u��!f�jg�w"��x��$p3���k����W(���O�j�%���E�!r�a��}�pF4��h�`���;�Z� t��
�9 ��C�A�E�����L���$S�h3N��b2�uJF/ ���VC��b�Oϲ��B��ݥ�(���4�����]�F[�!�\��n���=")'5��0o�Ѽ$x�H���nj�~i�U�⋓���k�R#����7`�!��d�S��p�����,���s�Y ǒ^��v%����RѮ�v��!1-��S���P�)"��^��Cȁ\�Z�d��PԄ+k碈Ml��n�>m�oH���]]d��QS@�A���I�bASmi�N�G���㏞ܻQWt��ta�E��TOTO2�H��"o����d�4��7�H�x�ǁ��� �_�����8qĽO�>�X�X�F��_F7;���keG�����k6q�=f����hɆ�f���Qo0}mK��v�c�+�#�����p����K����!��I�&�dC-�r�8w'G�q�����(��dzb.�OC����zN�>��?��m�a &�4���P0QȖD�cp�JW�"Y�\;��a�h���^��J ���G).���¯��W�^qJ�� S��fH��سJ�r�-��x��� ��0	���iiFq�ț,���Ǖ�_��`,�ށ �I�ON��0e���A�v�B+8���xȏ�X�Ua�Ы����|�A�ڣěN!am���: ��ŶKevΩv�#�)*i�A�����I��*�;�$ǃ�� �w�&��"Rmv�Q>07܂��vnK����l��%�i"�b���o�HmL�,8r/+Zr9º���cO}��T��!^��>���$��L�����$u�>�a��|
����塚v�G�738��v�q���������%h�M�&�7]�;|Y�z �g�}AY�՗i2}�3��X�ꕱ���0=�զ�����F�7`����:9a#%-����b�l��"�|�t�:���{&M�r,�4c�^�36����?GBK�L�jap��<7j���E@��C��$�D��샫d�w7�x�򒬡$yYc�r/�g ����շ�n~�XM�f��j�g|�ވ�<g�O(G�y�5h�o�	't�
6�<g����E�z�g��X��?��,�F}��0���\PϮ�sڡ�*�$a��{lY�If�X+��p�}b��i��0��F���/�{��2>F&Z�BB���t�F��;��^$�`Չe$�u
�a�O�1s�WO�:R�1�"���M-�8��x8K�z�q��4? leB��)��m��п��k,1�wD�R:D��EBJ)˧��x^��Nq ���O��[~j������f�c �pu�SGU
Fp���s"��UH~#Y:�����@|JJ�W�_� ���P`8��3�T��jG�!��L��;Χ5�෧Bj��!��rm�h���}=�Fb�744��x_{��Zo�>�A�xE��N���5�p����Gҿz�|��T C~/ª_�G���!�����a��2zdMrv�l�]/y��#���#9��6�-+_�Z�����n��%�`>Zh�.DO�|$QO�w|7���ϙ>��\Mv������V��}�@��} +x��,�<?-L2z�qҒ�9����vk�$�b'��;��OiIC��]Çt�����Ėd�c�Wv��������C�<\n84BKD��f����"���*�+O'�?qAr5a�P�7����1��ğ4�W��(Ӻ�+�C���\��HC��%î���k��n
R֔���x�rgX�sd�l�@8 7QK�Vfٴ���-�8�Z��d�_š�Y&��I��xƼ��mw�zr7����2�J�^��1R��GѪ��;�v�������l��.�mc�Ӗj%78W5Q����w+?�~֊��|v�e �`�>h�^-َ�k%�T�_�{`�!+g/�OמX8葚$}�Ϫ�{4���;�P�-|y�:_a�/=U�w�n�r�<�g]�ک/n� �aZ|η�UQ�;Ŀ��_�r���w�-t�����rhVxA����ť�#����<�<)�	I.m���I.�ȶ�	�
����u@������~���y��2�G9�*2��|�n��hy��'H+p����Փ�;]!-F\ �]�j�ZJ���+ʁ����di�����uB�ݝ�te�{��MZ�\QN�e�2S(yQ" E���gG <�O>{���B��f���u����V�[Y�9w�sH�pX�#��Y~P8F�8���׆;g,���#26������lf��Y���p�H�J��[��pǴV�Eg#��.������T���VҞ����>o�K`�2��UOB�zW�t���ޱ��1v�NI��i}��,��A%m�!�o: 
F#@�~�4r&ۨ7n	��=͍�v�Ȱ"�� ������
26��j�-���]J;P�`�B]�w@²e��ӽ��k� �H���X{�g�m��_;�O�d��U�ɭ~ �e!n�b�l���:���Tn�o�~ˉ;Wg381�Ã#b%�w�'��7S]��gg�x|�CO[![�y�:)p\�_jKq\���*��+};��y�!M��5g�3w�����;�V����=<��9�B��]���_P�R`F-#����d]Ry�����3�O�C�x]�����F�����`v�h���R��"F�0*�36|C��BJSQ�i]�!`klh���*����P��5i C��\�6��k���b*��|J�Q`<�����V�X�%�0�socQ�j���α� 7fUa��>3�H55|���2*�<�m�sb���ƛ�[�s�μ 7�JEm2�HQy�x�;F��=.�Kg����n+J��?�@�d�u��G5aԢH+k�Ƨʘ-�} ������!i$Nr����g��&�{X�siv�;I&=xhB��� #w�����af��B>a��g��((�48���s�>�yjz+|���-mѥ��ʫ����9��z����Ơ6eQ��,m*�96��M1��^�;��^���E������T�SO�Qde|����ga ��W���m�� V��hB��F�������d���3ڛV��5��OL��n�0� *C��8B����>���z��Yc���ʑ3�<|�x^�3(�\�"�)�g��%E��F_	N��^X���%
��� J��E���d��T��
�BǙ�$��fS����"�hAZ�-E����w����!!�gD�ea�%:�=�3��΃Zy�{��$H<�[���5ck�W��tH�붍����0ܓ���(�Z�˹���x�M�EO�UJ�~�D���^ �v�����*l9bnjp�T��U��"1A j|��2^oQ�̱S~P�\<D$�B(����i�bx��"��,��^������Z�5��s i*F4�Q~�o��Za���0R�����l�<�	f�v$�����H	�rr�5k�^L��x=mH����0�o��v��F6}w'�%�l���# w֬� M�V�;�`�;-m�hov��J�"۬ ��ћ)�"�R]����X"���������X#/�ڒ� ��~m�)���mq�-�3X �2��K%���
�[.�Jx���\M%�W��N1(Ǧ����Y�u��R 
��#	��qZ٧��!�	.;�A��@��M��3��YZ^L��-���X�aI��=5��l� �&���^�hz���Ֆ�썥~�t��c.r�((���wN�[5����,ۋ/��������<>���^��$�����61����c0���uB�"�´p2w�mR��Oq�3eP�N}6����f�M
����6�d��F��u<[-��8}?�[�&�<�0pq�*� �^�ʊ؏�hW�	��	��T!���
iЊ� Q���<�ku�<���X~�фD�;f�p�O���r�����N���C��?�Pȯ���}��U�L��ȺM�(S+���iN��y���l��&}z潃�Uq���=���g$J�<����BǇ;:���x���c��2���&��rlg|G�Sq�/��5���շb��9W"٦8�3?� �����UH/��8�[
p�D�u	J�)���k�e�Wuߊ��@f\_D)��t�dO�"s��i����$Kh &�)�������%KVx�@.�Q��^���<��	i�B>�U��a&��
�`���2H��<�����*(�)��$ nʩ�ڽ��
�WC���Fc�ƹ�Vo�<�eb��w�F:4$jw���Zl�ݪ2�k�B*B�	$��?h��Ԝ`M�|�SPsΘf	ݱD�uL��s2~�����[{�OLU'qܝ�܇�1^ڭ��K[j7��ܩ�oҼR�!}4�3I�xM�pA���Bb�-�⡂'��'�-V��4D+����	��Q&����#�m���efZ��}�>5{R�}ɀ��Hb�)�J�Rs��[�V��C�t����j�O���o�揧	j.��{a66��)sG3�7�T�H%����V���W��(�e�i���D��`�89��{_�][8f|�
�%ޡS��-��0o"��0��>�W�T�ip��5Sl�<��Pw��~��^�Uu�����'�;�\'�	�ѯL42(39D�]�qGѥ�v2mmc�MAV}b	��e��;CO6�d���?�
Yw�G�7��!K�u�B���g��=b/S�m�\�1�ۂ�X=d۾�l8zZ�f*�NF �$�Ѹ��Z��΂ƨD��e?��X���@eN�w��ov�5Kx�z�usF��WvŊ����%KܗU�����
���b���؉�%����~���r�3qj�91mc����UR��
Y'��w�E�m��ڋ�F��@��bӟ�(�͙�/���C��>���%�9D�K��@�eB�CXLٳ|����QY��9��f��V���({��pG\T"�d����I_p�E3��V}�Z����Ȟ�_.ޑ�U���2�6)�
�E]� TXiZj��Fg��o�J��4�W�×@�g�N��}�`�Uo�ho:��E�K�mEw�#:�k�E��s�i���$�Ʒ>\w����-쏷�����e��8/_�:���ޅƀ�1�RsJ��A/|�C�9h�9����uu7������Bth�Δ�#7���cCئ&xho��3�8�]�l��N��_c���-~{T9�;WE\�h�v����t9ypB��
� �[,��u�:��|�s��E/���U�?���k�Ր���k�M.����"kq���n����޴h6?wv��2.�lb�r�`~�"ʃ�Dg�a��q1�R�'IHb���i(��1�,�������i]z���;$��n0U�[��u��{��TO�����t0�ӹ�}�;�C���z�*�B�u���/��*#���S��/ah����]}��?ZV�9y%4�$	:2���k����������e�^V��m �����\�x�>�!����7�LůJ`k�P�8bk�$P "�6�������fh��,%�t��#��mF�����ܸ���]a(�;qP�U�����	sC����p����r�HI����w�(4|j?��c�g�B��-�=lƘ�;.I~���C���N����g��/����6���;�'�6��W%Qi+����Z��f���IQ�A��2W�-��z��s�|�E�{[�2��[����u���A�'?.}AkRJž�C�8���č{Dok�Z5�I)�
6��ͦZ2�_.�̗��i�*��@8%['�೨!ƾl:����' l/{�F�^-	���b��j�ǥr�y�>A��y����r�ш��y��f�����%b5^��x��V��؇����!�A�@�������٦�2�2ْmD�,���汹�ᖜ>�	 "�,�:H0z�ux	�}�����Qk	�Þ,ku�z��aԻ�!���o�B��-�,�U����E��`Ч�N�����磗���U��l!����Ǟ�����0H�+�g��F�4r!�<r_�$=T�A¢	vj0�CF�<b�E��<[(_�a,+�D�j�	�9dUo�)�c���:5D���;���8l�,ZB����;��$�)�6e���L��}�?S�ґ�!���q�{�UB��^�&�����XMt!THF*r���q,�:Y�WXN�o6��}7��c�c	\If�݉��h��ь��t��.��:}��1N�s	���Z��v�@b�|�G�E���Y�����0~�����V���͐�xA"��:�H�2�X-�,�Q]���W�m��"�$���0���ۦr������)��9��U�� ��jT����:"�`.� ����,eZ(�
1���Z�F�څ��gP/�R�)�{�E�3K39_(w�FR�� ��xgv�D�FzO�����B�k�j�=��2����dԦ��{�f����8�#�cge�{ճ�by@j�3����)�����2QG��4{�ә���_���p&�.��H &�{"�1��¾�&*��4�������bTKD��8>�o���:-����R�s~JR��`�6�3���[���|6[7?�v��6.·p���� ��8L�o��ڞ�8���&��d�m-�:�FO^#���y��������f��h2%�����4O� E3�S�h��l��#�K�ߟ\��,x_��[��n-��I�9�x��D�hat�8L��㷟S���x�/�׽�֖6��C�3��zE6<��T�TB��%����M�4���X9���?�߯k�[�Cg�S�J�r�֠�n��Yu��/�e���p���hO!���	t=�.�dDT��I���B"�2`�cS�P9 0zQ�'R��t�c����3ysHjEA�o=�G""«�*��$Sf(�:�oM'��:��)A�I�_>㱸����;�0tDW������{P#�q�T��uށܺ��h���Ex*�!�d�:���7�*�}��V@V�賈xi����y@�kz�P��5V��s��Xeɋd�oX4����8��?
�u&I�Z%��&���~��5lq*�q}�n�3��P��
�7��M'��ȋ�H�b���K�I�(���Զ;�����z���a��������`
���fT|��+Tio�S��c)`�Uإ�Y�Uj�Xs��h�Zi�|�u����4��{��P��"(����7�=��*%�~�����8��<�7��)#��$L�:P��hƫ/S���` Y?��t��mh�E�H�s�H�������
��	,}� �B��G*.Gk�p�h�Y�Z��Ϧ����,��C,Q�m0!3><���u�j	�hC�L�����èR1aY�UQ�d
:��` ����NE���~������L�n���`���[�<�$R�<��00_t��M�"�]��M{�9�ǨN%:��b��#^�lvլ	I��_q7��Jy�վa`��.�$�2#{�8p����:�M�$�����w���0I8P@���&<�x�`��!EM�4h��kd4�ٌ>}�d����EZH��\�1��͛_e�h�S>���8S��RWD0w��<���^���d:�-6|���6<��4>��Q�sn�1-��AP�v���|@�Ô-1�;>�05�,����_���f��N�(��B��0J1ƫ������>2ߵ]�ς\	��KZ��|�P�߻L�F�_?����O�~zR����D�6�ݩ��J�f�������>=�$�`���Eu��5�|��jc���;W�/A��4MY���?F)��k=�<gW+kV!�)���Gp-�g�Vq�.(�l*��z�o2^�8��1Oe����0$%3��ˮ2��*JC�.�y�f��9M1���~���چ�6�2���~),ԑ[Bɫ�˖�@o�����rU?Fc�� �sZ�"���?�ɑ_(����=���y�$d/Iŉ:�d���Be�!��Zb�w9"�Gd@��!����xm$IP{�XP�9���4��R���_ ׃�����q`kh�\�v72�q ���)N"㮌�v�E8(��n�p���Jf��Sr<jE�x�J���R����PBd�S����/�����91�^
�_�H��r���Skg@1���\�2�?�GcA������>1�ۃj�5�j�E���<�Db�ئ�`�3!|�+��Cw� ?6�P�Afΐ�#�F�j�j���_�-D��(�xA��;;gf4�y`�dƷ0=�� �c!ֱ��]�4$w=]�<��/I,���*%�W�W��^�s�'�}j�9LDU����f:ʒ�2��v�L�.�����(�~�4Z��_��YZ��*Q�⑊X��
YO&�,�jض�l�������]��c�6%���ߗ��k�;�fpG[:�BnA��&L��8��vrn��ᯫ�y;�.ַT�H����A���>���jL�&����j)J��\��U���_W	S��2���ϡں6�t�F������ϡ�O�a,g
J��Lĩ���'Q/�&Wzx4?������:^��L![�� �cZt~�����H ��������C�LlAu��ie� �#���bb���������~g�������ɩ����Βr�S ;��d�D��!z%����Mw��s�7i�ŋ��1ˌ�_hŎ|����iVmd�ސ���;eب���J;�]r���K��}�6�5�q������'h,W���?�pr&��C�
�q
�����yĕ�)f�C�و�Z�����J���:�Ba�ҩ'��S��xw~���Xu����j��6=!P��H���C� 49i�57NRG�1�B�%H�@}<鯗�u�?��܋��2������"��rH�E!�"w:���ٵ�Iz��s�<Q���"Ֆ�O-gv�s ��s�H8E��o��g�'�I��"	a�j��A�ʹ�����DK�p����*�1|)п��l��A��;H�˗�G����q��h�I�,��p>�X�Z�;4�r-��dQT�" 4w$�4,���&��a0}��&i��JR#�Ԏ��i�=�=alq��|���'9 ���ض�s��~KG�nR�o�؏������ Sև�T�Fp��j���I�5�h/���U�3�P�>��Jb��Q()��g6\��6�~��]::_����d�Γ+�*��MV`N�ig�<b�	}X���T��6�����\s^l��}-�]�x&�]��a㪫����zy�u�ߺ��}-��!o����b�c�zU&I�͏�B�u���f��P[���l>ޞ'���r���&����e=���r�����1ݬ[Cɬ�|�E�?�r�h>���f�r
&��fj�:�7� �wF�̈́��f�G��P������3VK�,��=r$y�m��Su�g��f�i͉hn3<	ȁn�	��I��aD�%�Kl�@]\�<~w��-��/ �f�n<���a�'Ty'��2���w�oyS*�	���&�5��2�ڜFaHT��Â�-!=h���j4�#N
�*��������,"�D���C���S��{�FI��g�%����f��e�a�I<��������D��������M����WJ&��w$�5�U�� ҝ�}(��2sR�:������M&�nj�5F��xi����t]ED���F �>�G�V��`���`d�|�
w@�G�fa4�֟��F��ttJ$��o� =ւ��ݹv�5X�$�=���P��>'R V�"SK/Ǆ{��WGǜ�
ϱ6�:�+�hU޹d��ݪ�ʊ	]Q��MvD�4�h�m���F��E��t��^�']�n!6��g�I�	#W~�8!�c����6���Okа:G�
�>����Q،�o��ֿk� �1ݤ	��'l�3ka�W���.���֡Q[u�}Ҥ�>�!�H7��F�2��
>/�~�w�
~�#t�8vx��(�[G�{)�^��-:��Y����J��e��)�R�S��M�" �/�w�¿x~'�7�Ά�>$?�p��+$�H���~��N�AbS��s���O8u�����2ϛ��zK2Ϫ��L�2���z)-��r��>�b;}����zS;���6N�V�v��5�5���d���;I
�����߿%�7�y�z�qGIӭ�֓n�~�zF��=_��B��L��J�'���m~����*�F�7�.��*��=7��a�J:Vi���GVg�
]e�J����i�����aZ�`)��1B�(�u�R>�S����X>�������K��{�7Ѭ�g�J�Y��}iK�:�/P���"7o�U^�^՚!4��\T�m��CI�vJa���x�z�6N��
ë���)ٟ
q���X�Q��g�	,A��W����&�99�*��*�G2�qi=��>�6/4�%6����u��&+�%  ]t�&d��Z��d����$3>��� 8��D���i�,�������H1��k��Β)zUA�X�ju�ȿ[9J�ub���@I����uX 5�0/^n��ۃ�?��dabL�/��U��܉����.;�/�8m�v�/#!���t(*QR]Զ��)���0~{=���⠖��<)��HD�����r�x�r2� ��;��V3u�Zo��!��`�$sRd�RS��<#�����(��t�ͳ�@�������-D�Q@�`������{���	fԖ����g�{���`��ld+��3��c���zU�3�����hkj3��XlxV64EB    b571    1ba0�Tsm������cv.*j��b�����Å[�|���5[ek��/ H�4��M7�'��l�?g�Qv�HM�"7����D�f���v~�_2X��C}�
l�$�WD�d���N������_�|Y����7����¨����'K��g����Bұ���ؓ�Ն�W�D��)(߬�TR�5��b�BX��G*8#�k���A�y����D)<�Bw!NW���Vһ?|]��b&~��q���=�B�E/�׎5��ϤI<�X�P��Xףj �R3��� c!(�42Aaµ��C}�y��"�ɾ�,�15i'A�y�K\Z��h5t_�4TH2�Qh�8���vLL)���E���4YPX������ϻn��/rr��R�;�딽�Pkd+�Ųo�l�g`N3���S"��_���i�m��:���4Z�:�e�#��Ҵ��oHr
�EԒ���^>�j�)���&e����j3�1щ]�����)���SXM]�S�t��L��Ji-9�у�*����|G丩��5ѭ@�#���&�]���Bm'��� R��;-�
����#׍�ez��w��W*h��������b犑�y�r����[2QjJ�\-�C�d77L����fqv��`�F���T� j�w~C�HoS��0a*��f�?����3jXV��(�aۍL���o������q��ץ~�������?48}�˟�eh� f��o~0z��� z��ǽ�S2��)�+r(g}��~j�V��B�ev��-�������%8��u��B7Z /w�)�c��K�T�����\.2K2���ο�J�+�Y������;�
��$H��x��)l>a������̏v�Z�q OM&H��Et_�l�EP��U<v��cQ��7D�rC��_��@�U��f�>�35����w�k����ϐ��+�"4�/R� 3EݨQ���V�}-��Y�<�z%s;�bBf��g�t��Jf  �����Y�3_�Ɔ��9�3����`T��
s8GFנ�
������@h	c<�@�V���e:.O�ڻ�yaQFk(PIJ��W��<Ok�M�[��p<��u�Xs ��l�5�~|���c��t�煮��|�����������wKh;��WY�t�d�"����x̔�4Ӷ"{��q�{!�xQ}O��e_t��(�n�.q3V0�A�ڐ'��uİ��'_��)֗����j�<H����TcTr�x��� ���jn�!;)����¸�	��r���@����hR�U���s��9^� ��\��h�P��@?9߆ Ow����4��z3yQڏ�ɷ�K:�st�"o6�ז�,_��fGΕ~���:>1�%"�~���i]��gx� ���.�w�j��Vۥ+8�� Q���;ax7��(��,z
�n��,�H�QK�I�`����I�	M3�����T�E�<Sy�uz�D���X����-�O1�;�-�a\�'� ���^Sb$�3��fa��7�M>k%X���/��[Su�w2��W�a2 \�#Y|)�TLi�o?��s|R��8lV�U_EQ�W��}���ˉ��Ϥn�I����H4���a1��o���u9 �$�!�]]��E��S|�8#�`2����\�
�g�^x��;4�ھI�S�my�{�^/�rC^�"�G����1�Z��/% �< -��_v\9��/B>ف�FY �:n�	 ����F�h�^�� �G=H6��W+�����wd Li�з���'WէK]�坘q�3�quͰ�J�ǚ�B�mx��TA�E�����'[����l"*����.�v�EnI'���Ǒ��/2��^��O64�5}5HE�U�i���
R[���=�洼�Z���R<��1�)2Y0���n��!)��}�!�y�,2���@���#��7rN��1¿Y׉Hݟ$7��I��f�8e��W#4�S�ݳ�F��%��'L��k
���2����z\��N�?��7�9�^��OZ%@�R"l�H�V��a�O8%C�� nX@��T̶R?TZ2pH�D*���t��`h,Ciճ�{e82Ԓ���Ns���x�Ԝ�W��IY��('�&7�UwuѼ��<���s�e\#��:��MPAp�l�S�>>��1���8V��o�%�܎�^閍�O��@���#�C�[g��� �`I�����/�����o��r�&���^����kCfB��8���BF��'YO��������>���`��0¼R� �^x��r��JԘq�.�<e�1�����#p���G�·%����nt`��|C��/_�}g�2�W��e(E�"�o�=J	r!�p?�e��U@��)��o�*~�[�;��,@%�\�-y������ ���o3�1����a�S�L�N���ЌX�OU
�j�x(�V�)�Q����f���U*�q��W� �X�Ȓ̭�JL=�*�!��\�1w�̰��QS��(�у�(h:�w�#:���\���A���ԅ���f���n � �RGgB��aj�G�Nk���|�Tu�K���i5�z��e���j`3�1�T�������Y�6dy�"�[~���i����?�Ȥj�.�����L�MN�i1����^@�O��ǌw)h�PC���5fYvu�Ͱ�2h�+�=��zj��>��9I["��U>���!��53��V�!��<h Ͱ*���3V��}�@��Q�K��`Y��#J#����,#s=mGr��Y���/����.���\��z�b4m�8�K��ue4�E��A��]�os�}``2��'zsۄ۟���4`L�<>����Y���b���O'��F_�9;{��A��g���l��,��/ō �0o�h���F �@�I�&DW��+��|="�o�3�3[��'�KI��PcwT��4�iś�I��2��*lX��D��#L�e��K�$��}�N�U��%ʇ>ĳ�?ڨ�l�9�@)��Z�	/��٣�oFMe�5�"�9�݊ι���7�W�D������D;� �{�̄��zvI��ؐ�����t�H�n�,�,ԅ��ݎ���e��.㕞��d�5�����T�#G�����:3�9d�� YcI@��ۄ��j̑��_��KO��q���x��3	�����6µ4���{,zPF�3L��o5���m*? ei1�<TIaZU^��WHR'Ì<�	���!�� ����
�,���b���M���q�~VK�^������K�^HG�_�r�p��G'C��k��-(���#,�QI�����&V�Uxh$o���A��7�>
EN���+�\JŹ����~�p���ڤl���~���}�4j�A��.�p&��X\�u�3TK�Kht #���Z\�ڙk0�vO�Tu��xd�.���y���x��je��,ܧk(�[d!�>GSh{�=�/ǽa�D�9]�K���^����_�}mJͲ��8A9���i�kqO��ӝ�JK�N�vy��!Lf��v"4������MD�r�FU\Y�H?��tŃv�WՏ�p�^�V�%�^v���#뮘��|ѥ+4'U���\;^��q�Po�r�Bl�%�v�g�%�]nG��k�����g�]*�^*��oQ�tx���ũ�.e���c2�&�����F"�f��my�ق��hl�ǵ�ly�V.{�3��]��!���s�s�:���� 2A�Z��#t����ޛd��l�_FxpW��I���B�X*�K"�O�욛�'c��㙳�T	�a<!�(��� ,z�Nd�|�"�Yf(��uW�׸݄#�u1�a#)UE���e��#W�Țݪ�I���Ż.m����;���x�� ���[��V:&��t�j�?4��.5�Vdh	ѓ�T���@l`F�f��Pg��3k�X9���X��澈̷	����Ć��Ĥ)��3�rs&f�jQb�U��o��.~�8EJ�i{���\9&��ﯮ��V'��z/��}�����4��<Ώ~<�\JRhĒn��r/Z�vo�������g��| ��y^A� �1t�׸����5>eƃ˭��	�l�k�\-�,�E|���ʕn���h'�Q���ex.A�R$��uR�ʪB
`��w]�j�DV��Wx��x�oPT�>6�5��#��Ek����hM<�N��A���@�����g�03�K��s���7�'�Xw�h�JX#v�"T��L�*VHyg�Іf"��a�l �e�W�,���?���%qx<bX���3�`Hpo��y%�����r��I
���H߁�����>-�q�y�2՘�c����אzY�f�¼10+�B��eFL�o���� ��?)�
���ظ�1�B�|$����@g���":����c��РyT%9
U&t鄌�ׅ��k�?�ԡ�b�R/t� �m�����L;:r�>��R<����%������
LO��@��4�'ב�#����
J�p;�����N�L3iЧ��u�GN���`���q9�1k��d��F~�z�Ev�PĚ��"�C3�I#�c�/D��&��e,s��6��yo�QMH:���mQp�2�����6��O�]ɰϙή�\��p���x����e|8W��&�!�|0�3=Õ����|�������Mao��+v�P�
,A,�����2i�f��ֽ���W�3l�����#T�^��8���a���Tp+��f䑜�9�y�TA�O��T3a*�л����f@H��W��4Y'��i��Pb�<k]�"�`�y�C���LcNy%Um
Nt��02�^Tkw7Ϡ��,>��G�Ya�oo��������(zyg�T���t~�N��׵������_���MB,CT�3��
��p�<�;��Kjm$w,XI��2 "�ʫ?�=4K�`���-��H�m�=�θ��{G?�H�p�;ױt`��F��^������@�ɹ (o�&��vd�����8��Ax�q�k�9��.��#Ȼ1�ӑ �i���k\���l2�_*�gJ;�)X�\A�d�U�m��ј���Z����*2�s�c��[ś�|��x��S�kY�Qo,���1@�o��%�}����i$ƶh�uxKI^	�@n��T;�󄣾ܽ�4���G��v;�H��&f����)��oF���m�U1�Dvˆޯ^?���>g���R �K�mA�i37œ����o�%X:��S��*�a�tCScd�.���b��N�Z�55�0-����;��j�c�	�a�mA�_����˸�A���Yu%FpbL�wr���L��5lJ�P������=��h��w�De�o9�5�v+d���̱+��ޟ��Y�[햛�a���ϳ�4��9#�P�<�ٕ���N#�^�F{鍸~��:�>\�����Z�׭����,��֡
�u���m����t��d o�V �J�Ҽ�F:�X��D�W���I8��~%��Aދ�ې	���@'x�3G~	_γ�bS��@�Wj�#:����V>U�ޖ@���Ee���L��Le��^������׼���3�>���kB�j�6�͔�]�vP|͝IA�v��0I�cz��_%Rw`�O����^o&)��#� ��͠9F��_]`nfb��9�FIOn�w9*�e���F���8@:mڰ�ɧ!pQ�7}�x`���2����g']�( �@�?�<�x���hT��o�1���CW��P#me�Fz�JM7,��?��_���^b��J�|2���p�Pw)��L]`@�]x0U�5���Ǿ��6���S�~�t�%�s�ZI�����̘�6B�N�,Ʉ&2��u����ݶ��F��;��ۋx����|q�Am�(��]MC�l��$R�(��|O��t!9%E�țj�q�"����h�V��/���g���y�Q�i`�v�0x�����r�v�Mu�`A�8	�W-�5�M�.�|=�_�V&���Z�͚Q5�RHr�񽆱O��f���ۮ3q�=��������(�rX�GOA;�JW�n(6��`� ��U�=���F�d� 4�ԫ�D,{�p�7]n�0#��!�U�A�>w�P������r̴�l��Xx1�#<�n�w�26+%.��gm�u$��Ó�������﫵�0Z�RR�N�v���濚�u��8 �2'�ǆ��l�ru����^Z��ޢ�����s�a%�%c�@??�^��@���ƙ���L�_{�e��:`)�~��6�2I���UX��!y~۟��'x_� D1F`x�C?�t�dі��_hǣU�Y	C�-�gx��+aJ��0��%�z5�Evl0bd�P�L�Ҽͨ�����r
��p9�:�__���gw�T��iE�̈́%$"��[�wZS	wZ������� p��3C�[/���d�՟6�����+M����i��"�	��g�Ȍ���Y�6�C���n|"�� (U���Q6���hU	���A7�!����P��IP �����)�#D��GM�Dh�|7�AB�����8mJ�K�$���cYI�Db]��4��<�~c7����Sz�U
�t}%��ך�~�� �F_�S�����޳^d���?5�h^򞖒�;�}u����#�t��H��k1oa��/�}9	Ǡ.��i_��5��\����qo�A�@8�����������n�w訂���|y��뾋���=s�g�!٨����^T����~�ͧ"%�I;O�p!���7��I�JB�0�0ѕ�����\�ۀ�6�bBR�O�cHu��3������f�yF'ްR������Μ�c���sqs�O�L6�3���W�.Q"�����u�����m(���,��,'��.�Yc$3�mʈlz�?������ �&�l:���Ŝcѩ�U��O���3*ҷg��S���X�>|	�qƯ�O��s��yl �ny �����#�
�������n�rq��^���R��@.>���| 1�Q�}j��