XlxV64EB    336b     cf0�T(X<ӣ���J@����OӾ���I9���I~��!r�-d�#`6J�?���G����¿M�:M�':f�S����(	^Mtuܔq��E�%�ǒK��B�f��o�x�P2�::��}�rT@AH�U� O��2�#"��1����Wd��˛��X����iy�,�s�-LD㼨ע	,��:�*뜁d�o�R|�:�/�q�.X�m�ނ���@�6.�����YH�lϭ'`��ogjB=��~�îz�x�<��>�d�Bua*D����2T��J4���<��~z�=7פ�bb0w�#�d��I�hYAܽ�@T#����c_�6Y+�,t����tmMP�@� �92μ1\�T�J&���a��k�6ӛ	��qI�R������ Ӄ�|U���R�9�~����/iZl�B
�5Jb��cC���64,����kB+���ͷ�4�1T��Tӧ�!LW0qUIa�L7A B�\6�:�&F�6���긵��yc������'#�ݫW�Z�r�Ej0��T_ߥ�r�!������\������?�Q����q224��Uv'���iC=�fM�6q)H��7X_߯n7��T��ϣ{��}�N��CR���C���|U��e�j��ʐ��VV�uZ��T�K���K��r�׋��&��Ӳ�~ze�'�J�Ҿq=���ޕ��`/UT=7�֖�2�5Y�)6-t�HD���e�_^#mU�jc�۳��Y��ˇ�����v@��_�Зb�;l��8��,��K#8!���4��K�
��E�~��0�=�?[��I�;��P���(�J����;���%x�#��X�{���}t�B�����5�ar�/��>�3S��k�������5��1������(P �V���L;85>e>�o���)�j�;=���R�����v!�R�j����{n\�+�8�*�JŪ�� ���S��TDA_*Q�:�Ib�֜�@�~l��PK>�ƷA�������_��������H�>��c�%�yj���JO�qy�H;d�AS�	,b�6M|� �����R�U��i�O8Qf�KI��m�Tq����@�Х�?�:��~m�dt3p4�1D��'SB���K�R�f�����u�K�d�����9��F/���G�	�2)3����	\n�Mp�8�0��%��b�6�E�sz�I��A�?�߶Z�����T��������JvSL����/u�%QXy�
�T�s��h�9���g2٦��zԛ|��H��f��;/t�+�B���eb'k�}���fE���4e��I����ߧ�𐊠��]JhL���v��������K������
���$
Y61k[�gv'�ɨs����'���G�&���S;�?*/Dx��Q��B Ѩ:*ˊ�'%�Y#���)�pP�PG��sy�L�1�����hF���8�5��L��:�9���Ws�6��H8u� :֗���I�'X��j�����b�H�Y�p/��Qu>�;C촻�0��CM�����;v��Xp���C�o��P?�n�'�,Iڀ&~q�\5a�[=����N���I[-Nܬ5�G>�Ǡ���ƹ�T�����ˏ�9:&!�|����-H�}�����:d�C�t��>����jŞ!Y���22��^��x��7�=YxR&��7��P��Tx�#��Zg&z�"���{ɷ���GZW���%}nTɚ҃���Vl��7%��	쟪:�}���,�F��O۲ԋ6@9�֟��&8V�c��.o�*�Sn�~ �̚��dE�a#C�l�k���x��ѯ�<���X}?�P��(�DY��y�4N~W�e�V��˙Ѹ��h��H-#���I�M[?N�;j)|�L��e�-��2}O*<t��G��<�V1���+R��k=LSD�<Y�a����8i�eMM:ՙ�Iɉ�P�[N a@5[��bJ5,�
0I�ure�֋��c�rn[�K��N�N3ޅ<�U��a#ծ
DMʹ�N_�<mX�M~�9X�$��h�P�ˇ^��ət����RY�!�
�ǖ��GQ�쩳p|6���K�����2�5Hft��QT���	�{����!KY�Oa��I�Z�g9�`������#�9�.UHx�K����D{�k�9�����s�]���(�l���� 8�g^�|�Tq�Z��y��H	d/�;��{8cՖ?���ZF	谏��6��?�d�� L�zբ�r��L¾�w��PD�����@�a��a~��(�|q�~����qp&3�G�J��
���ה^\L��q�`�ac7�XD�&��{|��٘�	1.V��S8�L]��P��_Ⱉ���~m�2��S�t�Jū���3�[������$���U�i��
�%��F� �3�}�r����1��D�f)*g�Mt���2�l۷�u����{��ݕ�"�Y��d�ɚ�h�$L�v�pTA��*�詔���Ǯ\��Bϔ������1 �w�#8�A���į)]��p� �	�����Qᑯ�e�=��b�3��xP��9L�m궀�|�:�H�t�9/�m{�D(��+����/���(z�w}���i0�F�_ǆ/N:k^.Sw���W�
�h�����E�8ș�)rz�uQǑ8mF���w�k��'�5� ���k����-ډ��Q0���q���5̛��Թ������ŗg�6U�h	�m�RJ[PkRwQ3e�P�t#,�e40S�]�+W��K��h��IkU,4Q ޿�P�uz�Y�댻,���Q�d�|�=�s��pIJ%2�����N�02��c1�r�p�T�(\��SBf��i?���&%�7�ֽ���Ac�����&�d�sǒ�%Kʃ�j��M��B:���DͯR
ޫpg�mj>:�Sc���x��;��ŤX9�c�Br����kpe}/"!��3�IhrOD�� ��kiտdth��~k�� {���Wk��ܟ��F��,~x|���E���R��$�=�!0������̟�	`�)�ї囓��������μ��OD\�����IBd����S����馱�@ع�tc fTIz9��,��k$1e���*�+�o ��C%	?�	F�&,����P��w��྽`�.'n+��`���g�;㶒��������'qɫ��K�|�7�7<GZH��,�@X��?r��CD�8}�w�^�\���J��D�oE�t��p���}1{by92s+gP��J������u}*�>4�K�џ�sP�4�V�MHF+:���