XlxV64EB    2d62     a80Qmcz.��5ΑW�:��eA��XVJ����A���2���NT�t���
c?�-ai��z)
P��+�i(霦j��״)$Db���&w��v�fy�����A��$&�4x
Y,�������	��x0b"=L�y����K��~F��?��_K4���P<�+;�51pAn����'����>&�4Fe2x�>��?*�'�:d ���m���r�L+����c(jTdRL����o���jO�I���n��H���h%�m
����y(,.�*��K�YHfZ��I�I��sŅ}#���c/��.����_����<���2d��2_
(����ז�ͱ���n7��fY�r���\�E3�{(!
֒�UW���5��NCS����q1��c�!�n5�ԑA!ji�ŵ:�/%�뾋ue�|�q���,*&�[��Y�����C[���:�"��X.N("}����Ġlݎ�H_i=I`�z��h�
�u�HhR�����������vdx���CV��S9����в�����1W
c,wfIz�Y]��R���C,0�U�g�����2�z���%�s�r:���++Տ��4�\'􈍓U	%�Qh��r��˚����,�O�o�����W�v�RF�C7+�D�ْ̖��LR%6p-e�#q���P�G����{ն��7)�b�7���I<ˉ �x7�3�}I�D����]YX����"
h�b*6�T
�Y����sxtAS3<?�/��9��X-v�X�S]v�������IF�T-Bv�V���\��ӮȢ@Q�!Eۑ�Y�t�F���*J�h�������u��d\D����9=>��  hY0FEՂ���ŝZ!^�-�x{�W��4`�y�S�䋵H��YN '��<
�E4ml;�$����y,�5��h�=��y����&���ܭ����H:i$0]�{f/��%��쉬�+�T�h�#���K9���E q�Z�_�����7�HFI�b7���u�N��9��ܳ�Uݭ��A\�5��і���.=��.�XB�AP�j�Y��5rL((����L�9y��b�T�WD�����B�щ��\�v[?����̅��[A�/������A?��U-<�u�tfRm�"��;������⼔3˟����-O��P��dٿ�A֞�M�8��	b\��le����>�Y����.0���m! Ǿj���o'�Y��$(	"��dB��Y�\I������
I����^^�e52|��EJ�w�|�A3s�2��s]����V+	-1-3
�F�.	��e�z
�D.8C=��~��s���v���-��}�w����D�Qs��
���s��ŸY�s�ǌW�1M�d�s�M0��lJs1%?W���";w�`�/�%ceƅn&j�LOyX���X������{cA��4�������㛠�m�;�r�{�'ب���Ф�v���hm����8��ۄ��+��H�����P5�d���l���TcW��u(�_9d��!�S	�V��_A04N23�i�G����0�< a�Q�ˀ\�����g��?���xJ��.��XN�����F�cu$�o3h���fز܋J���O:���B��i/�N�,F�C�Kz���ٝQ�g�����˖�V!2xM�D�6���@}��%.�y��Ğ^ĀEo���(dА<,�e�"�F$��K���~��:��v��I� �NT�#GU��+Hl5W㭯ᆊ�f>������	;c���@��|��6U1�˦���ѫ�c2�f�&}k����5�j�ӧ�b���^�י����o��^�rl�&���	w�y��47�t�zJF�zHJ��R!�����6�0Z���	�STܮE�|j�<��Q��l�`)q�"��)A�[S���Ga�"�;��z�{�L�Aн��T�S���~���H^�u��g<%MvRu(/����J[�0�t����{܈@Q7��W�9��`n w��b�����A�g[�����D��=X���$��cPNWN�Z���u�
�{W���y��M�����c�6i3���2
W@�29��nH���E����"ď�V(���Laکjle��|7�,�J>�Ä���빫�H�c��]n����>k ���CX�M�R����%��P��R�R�
`�>����;:i�9 K�XqxQ���69Ӕv��c�DR]&O@����?k���1M���4���?<��K�Tn1���!���$���u��J��x���|-l�3!n:�LB���՞w/�:Js�'�"�F�k���Z�8
�dp���M5P.g,}�p^�C�Y��݉���?{��&��]p��(�� ��c���?Ce+�M������&���VEd�W���Pǔ������	�(8);B��G|�R*6��vU�SI�/��B$�K�b
H#	���%h�����&�@�N����6�|�O0�<�a�A���(��`���La����"J�,��IP��\���Xލ���g笢�����NG��������V�_1����0}�h��忛{1~b��}�GPJ&�j��ˑj�݃���B����rǚu���B�U$і�"���U �+�v� �\��n/P��