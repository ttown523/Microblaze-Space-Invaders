XlxV64EB    1e41     a90d��°̖�ߧ�G#D7�����~�kfC��v	s)ͳT��G*h<�}J[
�(Yh?>�2n��Ǣ�������tw�D�w���)#$�k���!O�+wx�긢�!�m���(�"��.ʥ^�R�!s�5�9Dзð�`"l�Ӯ�w�oW��x��c�MvN�A�1�50Պ�~�fT��C�:q0"�}RU�=�FN��P���ʷ��m�w˫��a�|ħ\\J���E_�4�O?����U�=���
����X/\+�/g���V��j-��*�D_�A(E���͚':�0H�͕S�	��h68�R�A��h��*L�,w)���傯l/H�yQRx��O�_=�2�����̯j6j���u>��g�P�������p/xp���Y�����a�2�{�iI���<��=�D`��1_���w�"ZE�>�j�6��xTw`���70	꽵��������.x@�[�9K��Ι�cp?�4I����Lȕf�1�X��7�'v�N�J����AS5FR�vw�ݷ�_�0���,���<O�e���$�)��O��L0�]��D��Dlde���V����ӵͤ�=F�)�P�,�#]& �]�������X��m_,�ư" �M�0o� GfS'��_ܦ��E8��`�g�1#�~� ��Sxnrv���˗Ε	C��ӡ�k�Y���_8��v�����7T�_�Mf��� �ov&� 7DG?ګ����O�^��h5��f�� 8��R�٧�ހ}BXk�����N!˒�9?�_T��juBɅ���Jcd���4(�D�j�K��N��:7�֠P#L��JL	�P���-&z7mƖ�-�ֽ͋��C��<&Qf��ZR6�IP��6��M�����\���¹�uG�c�=dFOp	�z��o�8��%~l�e%_[	"���G(c��+T��u�V�LPk&���������0X�8�O4�5�2��b�j&+y�Ce��.t�3����[M5}��� ��c����=��$f@�7������)�K�v��:�2Pҁx�5�)<�ջ�x[���f�ZS�YP���|�X9��X�OI��ֈ��p�s���`13�j�A�j�yE�O�lS~���0����U���oz\eK�O��Ogõ����#yn.�,a��_>j�rAC�.{������I���r�b��<����8D$�Ss�Y9���n^I��}�8Q}OxY�d��Դ���X�['��:B�|y�ŕ"p	��r�pQ{M$��j�p�>Ӷ��AkBt�C����]t.�i {�gC�q�&�H@p�z�TހA���Z����^s:h���F�m��b�q;�Q��? �z��[�`�u�d}3h��)�&�tZ�>�>A�֋yѨ\����I�1�����H��-ɦ�bXDw�Mc���+IfQ��^��<��V�xRq�锓5���m^5��W��L6��h��030&�߱&�!�а84�����E/wp��L��sT����[7��:��I�44X��!䇆a��_L
Xŋ�'w����i�"(N��z�QOb!�-�e6�l`���B�& &|�9ީ)��̀K�k��r�M`�-�fk&�ܴ��$g��DR��Ma�3l<q��� ^OtO"`���*jA��-�����+"Y]w�_��%���$P��!K�:|̗�ҶX�u�L> ���ӓ㞹T�Dg�O������龶���/��Z`2�S���ޘ{�,��O�_�]ѝ��T�G���6�1y��Q�8zZh3"���rv �6�Y��Ϋ�M�R����a|�{EO磱���/�_����zM^�(Z��ή��V�қ�Rm���t�a��fkl�q�QcS�/����ȻF[���Q��nWA�ž���8�x|Ô���!���{�'g̺�6�y7�K����c'x�4�!P�ހ����c1�-L�Y�)S���|WY�n)��y�Y���R����k�M����J*���������n:�{ȄK7�E'e����1+F��7Z��^YaM��������*�'� SI�������)�ίG�R+�a-�PM$��kC#���3�o,CI�Y�?ݝ.�LTD�.�'U$,��峖C;��Ч$�X�-����n����?��x�zB+�hA�S��ĕ�D�LF��w��Jʅ�z�jo��a!;���N��Z�r�PȾ�/�<��e��Ԓ�+ל�xO(`(��{	�&�`���"r�
�j ��-9}^d$ͪ���c�"���\�.�j@6z�/�Nt��!nr��T4�k�KH_@������I�I�Hے������/�D=�+V�~	A]��u$�yN�0[L���YG��[��������{/���cO�緘��?�H0��^ E"<��ϐ* �Da�A�S=��%�G��9
��_t��Cf;��r�����{У܌���k���98��9U�p�`P��]؏3�ۡ�(�4��_K d{5��&��]ͥ�����7�y��;q��{�v��S�>3����ff\^������ M�9N ���m����Ѐ�*L�-��sL��4d� |ӽ��Â?���M#>43��} �r��*��i�t��r�兾�����V��~�C������Һ��3��_�_� ���VV��p��̤XłV�/��s