XlxV64EB    8237    1480��N"�KZ+X��R��$}��SE-�
�#�l$�S��f��%�A�޿l��Żv���G([/3~4?3���\���x���Sp#�X��[�&ǒRK�~d��|g��tW�N`��m��FO�ۅG����v�o|�Ԓ�>,�ծ��x���br:��IId��K��-�'< �5!�!���ʍrY/��p@�b��)c_r�L*�5V�u'�g��E�D��e�Uu)�ƚC:9�q�|��%�r��� h瘄�l��{L��I���$�$�}M�I!�&TW�s��!���k[>im�X��j1��a��q��Z��A�uZ�Y�E��Z�S�h��uo�M@Hg�q��#���S_�4��>��S0�e�w���`�D0д���`�6����r�y@�YT
>י�b�{��_�������q"uL��{g-R&�ph�k�8��a5_��EK'�>�/k����Y�Y�V����i%#��i�g{��NZ�(��gp@Ƥ��ec>�ci�q������:=5�F,��cc�)9*Gg�ь��ܗMb[����
V���y�&�w�b��,���q��\p
�@;H�w#�$m&=��b�N2qh4sn.��Nt�#c��t�WBsp��_��K��}U'�ʚ�\|L��U�kl5���wx-7Iy]5���_��r�ڻ�,��Ϩ�Ȃ��d�5+JB��9�K��<xK�]E1ٯF#閂F��Q��n���/�2S�d�SW��d��p|������ݑB���!Cl�`n�y�f�@s����!)�h�Lc�;zQW")�KE�g1�C6GF�4M�⤚�lt�Kb\ײ�DC�Y
�.�.٫��FB�_�;FáNd�ck��zF���*�V,?�7�J8�<�<yn���۫9aU����u��S3�<@����\�̄؋r�>+��%�����=( *�< x_�kwh���3��x��Y���,�J�i/�C�(!��yV9����!>�K~��ru��En�o�r��OS�
�7���"�1v�Ka/$�N;���mW)��G:��O(\��<�I��M~��~v��?���؋�X)�Y�zn{?M�ޥ�8e���&;uO�ү�2�M�p���"$�ɝ����;L(�q���N��l�y���G�70�#o�b�n�mZ7�yi���-����p�q�k����������T�o����g�����,}�y�[��yZ�%�&S���C�v������KPn@`~g�Sϸuh����z5#����O,ԓG����,�H�5ͳ�w�6emjCu�� +K,,�+KM�ײ[);7/��s��7p�~��V�iF}j��������>QwlK��y���Uz��>%ۙ�G�2�'al��k�`�c#�:�y��;4�ڶU�����~؁beq��+���a��\]"7p�[v��{k�~����>�<_��ME���|���v��_
�*��\ll&k��*MY��
�_��?��φ�y ( ֚s�e"VEC�).� >��lƉ������P�t�U*I�~����l�R\��Z��
 �&S"v�#:&	�J�u^Rq*���!Q<� ���gy�Z�dg<�!ۧϞ����cH`���5�7����n�aD�tЅ�nP7���W��;b�������	��Pi^�_�s�xێI
�n9�=-*��'�V��=f�5#:;��j`Q2�|��^��U�f�W&�AXy������.���}}~SW���i�E�uN��d��g�A�|��;��Z�9���oғ����}�ܴ�e6��};2V�XE����޴r�*������F[�r��e�`RC� 4�rb�;�h��Ӱ�NLM2Q�S��L> �`uBړh��b^V������AMn�^��
1d����[R�=Ed�n�1k��� ݑ�S~��XW�D�J�k�@��"EGE��4"!��������xj����ޏ�W��������C1v����%o�ǖ���VC�Bk���}��Og��$����W}�3�S��O�P���K7b`�ima��.�f���cw�y3^��w@-�Mߣ�m��F���3��ˈ=�5e&7�(�]�-	�zh�|r��@h�+_�0b.��k����	�����D4���k��`�7Pɷ���WA7�#+�Gyq�̣zO'�(�wԨ�W�y[�[��`eB�)��b����Y�þ
qB��KdEf^�/R|�K!�-,��`��ft>F'�s���yX�7D΋ץ3u:-������,�ـ��q8E������Km���x�G�Xˍ�B^;N=l��EB'�0(,օ��왮�ܖ��Z�����+�8C��X��pa�N_��0�K)�)����o���h�c)
]=^�рfI)���щ�+�� ���>��!.!�;^7��E.��)�}!]�6��9_9'D`��[�����̏LV���;���?�P����[!^�1�b̙~�|1K1ߌ����҂�vLf2�N
\"SP�V�zn,��v� ��Ήվ��w��V�1��E��|�Ko���Vv��`���ȷ^f:�g�>M����,B'1?c8~_m-m�,ܟ����A�	��t.�?+hW�-z���?�UH;�CF%��k;����5}2�S��
���n�A?�p�t���{4:��K��2F�:�7�_`!*d<�b�Oab�5�@��l>Hs5�8NE��U����̺DR]�: �Rl*y��|ŮG�UJ6kv����_3�K8����gd��l�#¼��|���*t$Y���1�u��*fuzyǕt����c�lۖX�I�k�%l�)�@�l�ȧk|�F��À�p�zB%�y4�� �H!y��
h<J5���(�G9�v�;uk�,|�u�h���[�f�oF�ՀW��� �>V�o̥�a��@�9��o��6?�'�ے��	��fݽ����\uzZ�Tgy��̼�䪲��PZLKf�e��g��L�O�@P,o�G��0���vF�`�Y��=�?�DJ�8@�R>�t9� �k/4�(T��1D?eݿ�H{Ż��#� L/Wp�����/�V���4�c���Wā���(%��$yu��*s�`��o��4	W^Ƿ2�C���r����Qբ�
���x�wsIi�����3����>(�����K�+�Z<�T���jEcs����!�n���m�iHx�H� �Y�E�8
#|�C؛$U��P��vRţ�!Þ{�]�j$��B�A�- ;$b�����[9<�+?8�[8| �ב�������x���ٸ�o$c�ʚl�\�V"�&y��KE����<zrC��ڗ����,�1ǯ �lzr�.� =�i%?�%�s;$�D�*�%�Jgb,��9�"�XM��M��4z.3Tؼ��1��\�`5�r�����\�Nz�D<G}�jt����Ǖ4�1����=V�/:�a�"�-��i�NE��
�I* k�u�	���P��r�+V���r�Wc�L9T8�ڪ�ƽ�ot:��x~1g�	��n5/#���*�#O�Y�G�B��7���08���n9l�����j	�EN��>#�'蝒Z=�������-ov-_�|G4~9y:����%$�����Y�>��P#N|�|t����Mb��@�;�J�G/n�%���2g}����R`T6���	�*��E�9����x����)^�E,q��8j�����N�W����l��,��ͻME���`���<��Z��∠�Կ�骾�hR݄!����IL��3	�o�Oux�ʻʾ�<6��DZF��{��t�X�Z�����JO;ݏ5:5W)�u����|��;��+SF��J�vx�'��P��e���v�S@�{՜O,X�;�����B�\�3d�X ���&�`�;�.�e5j��ѥ��e�8"�Z��=��D�mF�Ø��4Da�[2�9���	�5NT��'�g���F�M����O+BNN�8�8�Jk���t��4�Ҁ,�)	�����(Ln{r�N>�ꖟ�uCK��_��ng�@��;����(��pq�5�cl�-C��(��|»z%qKν{<�l�F�����g�!�.��&�KE����s��y���ѶS��}�쁒i�/�_jLS����n�E��j��<Y�ٯ�FO����������B)Ș�<0H�xC����]'��:��=�?QSn�\��"{8UW�r��gu���n����벏��I�ʌd�2 ���vW����^��=Vvk�B�V���R=B��ڈ��W���2O��r���+2J� U�R�Z�J�+�������$��.S��b��{�=�œT�ݧ��>�SN�|�����Q�
��^�� ���\�?�~�ܬu
Z�9
��Ξ$L3��C_�d��ta�\_ !F�(%\G��i�UZaђ�*���h7s�
;��BZ(�n{N��`F�<rw�9�G��	J��.1I�� �${��*��W0s�X�)ڸ�RZ`ӎk��ʘ�S���&X���t|]��	s?
� U4�2��h[d7Qއ� ��,�
�m�����*e�.q�k�ED���C�"���i�c dҴ���Ep���Nw��>����{#������K1g����G
s��0rpIK�$_��E�X3bƷS���r�7������>�v'�b.xy�	A��ݘ���-o�m��;�\i�]W��0|�v�����0��}�6�F-�}��ܺ����=��y�=�D������ZCme\�lw��u�(9��{A�Cʥ�����<��^�R���+`E����o�8~m��iK�s�w���?B�D�B��#*��n9��zR�+¿(��V���,8lpL"�{#��E�I͡|���Z.����O�~]B���%���=��s&���և��f��W�i�W���~��64ު��4w�s�\�I`?�%���Ɓ1�ѱQ�D���Cv�82�֤7�s�w�b��vm����?�v{��*�{��Hѳc�O���n*S�?H4��F$|cc��%��R�Y�V��AkR���L�'>��U��۩ڔ�Z�;8#d'�A.]�*Wy���A���ě�0j���Z�i@86E�g�7��,����1Mw=�7+��bA������`㹁�ɷwH���eq^ܦ��շ��,��M�S�UJ'�;ם�@r�G��G�V�λ4?�