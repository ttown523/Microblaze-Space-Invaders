XlxV64EB    18cc     8f01(q4ɢ�Z$#�=ʡl8˾���4>ʬ*f[Icnt�f��`D^����WC5�U�v�[�*�̂AԒ�|\�)l#�� 9=�=0v���2dy�y01��7S� �f8D�w��e����-)�e��n+����;�$��=��$E�1E�4�}Y�Z�Nȹ�0I��'hO�G��m%�0AL�q�����o���������2=DE��Դ��9&
�5�ok�S* 妅��d�r����((U��=��*��]Ǣ}Mu����n��w�w{A�u�C��j{/i��$�W3ב8-�b���s%��d�fxT�8����;�c��ْ:����|��+��@/��Ӿ=��G���3d��s�K�B���--1ϜQ,��R�?�K���#06���Z`�� l�~���sn)����S��!��!���K��I�z��=�_3��qQ�^���j�{��@��t�c��{�VM��
|�b�߱oo��Ak��\��g�+1���܎g�B�9%6d�V٥0�-�	���/
TD��>u��,@��"5�&5���A��XODLfjT�n��'��Ȇ�}�c)ug����7�V���J�|܆_@Y\@��� �Jm;1yJ(��G'�w�d��T��OQΦ;��H.���<}8�r��e�?П�+>w$d���Mg[�v`Lʃ9a��a��s��m�w]фx�1�����J�h�L�E��t�ȁ�ɝk��K�O�J�tm���R4/�[�o�J/�ƴL}b�>T2 هF������,a�+�/��J��03����R��+�����4˂�����讻mj<}xg��o5|��T	2�>x�e#��c�H�5�gh���W��������&H%��e*kF�#zN6�5R��n��
��ʿ���r�C����T��J\�(���@���}.����{�2�����u5&~@o}�8�S��C��_յ��xct虚��o��݋��d/S
ۢ�[SA�g��ЏhH����Ɖ�c;��K����]�i���d�o`99&^?V���2j�k2=���QfT���'�=xW�%r͟O�/���'�O���o���s�;�BS��O}��ڜ��4�׷G�+��0�eO>�x�.X�=O?*aƍ'�!3�p@y�v؞5�7_�.��U,�s�l�l�9���j�a����5����i���G:g�-�᪔k�zs{B�eU��9��Y�Cb�M6����H�1�����as/%p�첱�V���Z92�_QkE"37�@.עx���^�ÿ��y������X��&y1X��y˱8	ܳ�%�h�ڝw���j�<.�w�u��}U�)f���a}�j����]���q�?�N��/��Ke���~U��y�����mI���_ѻd���o"�`�:V"�	����.W-O�����w;�r����3�� �q-��&V�e���B���d-��MC�$e΂�E59�z��om�$�$DU]��4�lp5�"s.��1VC�q5(�z�{�!�k��35'c�_�!3p��4dF�%d�&e#*'ⳣ��9LPu�:�*(�B�T�?9[�W��� \�e�=�����0d��$5<,��ݑ�鉿����
u�8QP���y���x��,Kș��Y�4	]Su΅D��D2�G�l 4���ZcP�������*�=�cĄ�����7]F^>��zG���dh/�CM��`�;S!G���w�Ҕ�;ֱ�*=��Ju��K��q��������������Db;�����v��v�|9�=�mɵ��V��)�o\�ι��J�SGg�`���Y��ia;
/����B�Ò)�<���m����&�L�["���z!����eS�V,��ȷ��֜�["��2N�����8"��p�
f^�Գ3/�,�Z�@��Հ�[?�qg[י�I{j��E�ɑX�ri��x�I���ԟ� �F�I=H�rX�w��s����ۜ����QFt��@~�`�&��zBO]�'��3�ȮfD�o��n��[7~�6�r5�q�2�-�4E��}�1\�KB/�-��f*�y�d>-��7���S)`�鄌Fk\QƬM[����ڟ�C]z�����ܫ9w�ȑ#T]Ǎ�%�y�<=����g$v䲞)EH;8��z��k8��/
PL
%�V�^�8m�V�
�=�.��4�;�����k=��в|k7����)tތs!g�������
�C�EX2mT�Y+�$���E����x�X@���8