XlxV64EB    26e2     ba0k���R�	�
���j�$�H4��vYܙ���#f��k��\��V{*���x�3=�v���h	���3��L�ê�ΨoȦ��E_�'���x���c���jv}'wo�#�B#`�L�<�Pu�?���������WZX�F8�b:قC�B�+s�ysI�&�l�9�=����r�J&�J�`�����v/�?�	8�P�T[l}/5��5�K��0�Q�C�]�C_��G|���7ac�9)��s&�_O�)=���
��x��Hɨ�R8���ZD�.f8`3u[T>�7}��3P�NE�ogRs���jht:,����|PC�����ke�g���0�-�ead#&�{�'�%gu"ۂ8FN�Q8F+1]��Ќ35��4��;V�it[��Z}1
0�#Q.A;`�!8j����Qq����4� ��u�{I�f�*�k^K���kJݮ�)q�����=���7
�L����׆=�^a�v���W��f�l�|�D}KT�7�]�u�Н�wXv˘+�r�����u��|_�M��(�9�����/��n�����ۘ��Ŷph����4u���G��f��R��+F'�����Eo`�fV��#N�60�90���g �m7����Ь��X�L��2�ZWw��@B�ķ��i�mamp��#�\� 0��9��z)B��B��l2	788����������8@MBI�ͯa��䈑bH㯔�>��s�S��^+s2�8`\<.z7g�w�����z��pJ�{�n��^[���4�J� .�Y.���O�N��G���i�v�y��y�p�������'3y�ҟ�D��龮�����J�D�Anݕ�֙����5c�(��-��v}���oV)��	��L�� ��J�v�� rm��x�w"�,$F:������	��}�b�:�oI'���o����.��8%���,���[H����2)��M��j��v�������.��������f��4�)a�y�?�ܢy�^�Aʞ�r(4A���l�匇�G�9�C�cZm�a�-�� �iH����!!	c	H��=��t>��%�9���5{O�O��:`��aa/���C}m���TI�
�Չ-x��"��J���������C��,W����\�	�X}��	Z��}��J���<�l�iz_T-�\���[�f�TE����|*���'G��:���	f���u��)9�����r-�`���c;θB]#�����י� �&����#yep���VF����N�v��N��
��̎��3����P`kO=�� �����X���;����tv�Bj`ڽD�}NG1	�b2������P��_V�v��P�PU�8�5�O�N��z��^��ڽM���Q��"���H�h�7�&�/����4�ࡷI:��Ă2Q�Ɠb�ئL�x#�n�]��q��lb.�C���O�B���1�ܢ]��a*�����V��I'��9y��W?p3O)\V��qK�)p��X֔8Q�"�݇�S2dC��Z��3�]��nҟ�P���BT�.�2�ϋX\}������*�Z���&��H�4�Ɉ���ښ]Y�4�뵎hwT1qX(��D�Eڨzve.����#���]x;�vsK}0��nI�/�b����:��Ϛ�m?2�Ѵd����o�S��אg+����p,KJ��m6|pn兘�����2�p	;�&o�yO�}�fs����
�<F��|P��y��h���S�j��{�܉�ᤡ�T�������\�à��i����?�tՋ��k��̽��娭���uk�f�!z.��)�jK2�p��y��M��g���6#wn|^{i��U,JY1�l�����[��F�x�Ӊ�݋Ӄ����%�3r �Lv�����:gʴ(���qY�૝����D��:x���9����;�B�e��5j2j7T�����761��0��o���Da���D:X��M��!=�t�м8>v�n]� �#�$�Q`��h/����1��|%��$_�u�6���TT���pw3w��7���p";���i��������%Q�p6g��`�x3N��=K�)��q����Z�p�Z� l�8�lz:�;�w��r\�Op>��܌��&���ߍ��t��q�L��e�|�LP����ٖ�e=���f�?ڏ�,�8�I:�QU�����W>Z0E{�v9��jb��<@��ݒ�g��g�G��_wBJ��Փ����׭��x�+M�N��|��j9_����I��6
��U���9`�C�#�����G�<ꗢm=�{e�R�����$��ԗK�R\�zFC�S�.�|�ٴ�������|�P�8��#���7�٣��yl^H�\��&�I�F�g���R�<g<�������X]�ݷ�!�q0L��,N����۵YГ�H�M�UG.��L熕����7L���-a_h,2��<BV���Pd(��e�:f��.�����^5�����n�:�A��	�BwN��N^P�i�����ݩ]�Q��v��6�\R���x��e��(���MB�\E3V��	�X�t�;�	���0���9:DS*�ӣ[�uz+0^/`��O[E�i�����~���4�ki��`�A�	���%�ߢ�<H9�t�Q���@�U9�ѻ����[��7��nA֜R)����쫔Du��Q�Ď�)6%�L�>�a�Gk�@C�A���~�z��rс'�@�S��NA+ۍ�W�oh�N�B��| �9'�^l*
g�Z�s��%J����]�QId^n��C\m�c�2�=���@bd
v��s��z�wJs����|�0�u���}�����smM*�Z�O^遉��<�n��X���@���YE�SI�A9
�sK����VTo���E�ArI��~�����������@Z,kn�F`3pU��?F.�._z��