XlxV64EB    5ac6    1280�W���>R���0�9��������Ȕ	��.{3�|{e�K`!�,����D�M��44����f��b+��fSw�3Q�7���:0}�8Y8�������=���v�g6r�|��2����"J;k{�R[R������� �Cٲ]+U
�3ϕ�~!��b�b���m	�S��I�Rzq��'�@pyF�h�&Hj�� =�6Ԝ!�I3�r����#�C��T/��:;�b>:�e������趗,���L�l��o	E�$*ӧ�lS~��ɽO�X��M��2g�P��mY��`<�e���BpQ�UC�^ifJ�W���K͓O(�2/PB��7��rY-�͑��u1Aj�[yYe������RI�\O��B�c�wzU��͕.�;����m���W��mnoYN �&����@�L�v+������6��I����y����8�4DO�][�?S9�"	t���_�Ԝ��n�'�8.�c�8̐߯��q�gq(ƿZ4V~�3����"~��$$7(h�b����;�i�%u�*(�����[YL��<�3m����uk<�S/�6�4YŹ7�Xos'X>��1jCU�_ڿ¬�I�-����	��U��w�����o��G��-��(JZ.����p�)���Y�������{w`�D��"ho����Y4�E�W_����>^���$p|nrL��u��j#�rl�t�+�yI:b����4G�~0��`y�[���7�xN�ᮾV|�k�"�D��ŕq	i� 36n�G
���/9Ĺ/��qgF�F>93q�GІ����>�.�Kk��+����=Oi��G���[�(��� s���bބ���q ����U�:�/*�ڿI�����W	�/.��1>c�����k�W
/O���W���|�|�xb�Nkҵ�^;Ȑ�$��|Fc�{�"c�ܭp$����T�q0�h�/I�-i�>����Kp�?40�g#LC��!$�F�%�i��1��ٚ��n9y�p	HϜ�UH�Z�&�x����)ɆuA�~�m�!�3c$(�(�e"��~�u� �m���Z?���J�s@�ߙ>_X`9+��Y2<݉Z�x��Ϥ�y�$p�H8F�P�,2�^\���7�3'O��z��	<g�ܜ���\�V�ߜC���J�o
)IJ���ds�W'C����:,fX�Et��[�Ԟh��9jՉe2n6��[�W�������ԍ��a�Z�?�D���n�����I?��R����՝tJ"
Q�s�qJ{��T&\3Uh�kC~�'/`:QD���COFv�r�*�=i�(�LH�D�:L�/v�>��]�6��|EF:WF�xI+R���i����F�w/��r��ոG�ߞp0�yH�*���<�:���<����T�1���Q��Q%ܘ��s�}f��}�S�T>�%`��e:�>���';�r��Ly��Y�Y�HD��G#��p��2^Z��@9��\b�d�/d��u��?x�#LX�i����B�H�e����Y;������D��!*�B|(�&�_�[L�:�p�����
���~)m|�~:1���.��lg'�"}ס���?�Ԧ��t���ϛ@�W=A���x��C���(?>���KzǺP��*A��Ox�n����%�+2�N��诳9g^�q�47�%�X�v�~���n� k�'I�Ybs��#��t��G��5X-�Li �m��i7�r��'O�lB,U��w~���8�2�s��T+mޗ4�k��\�TI$� /����WI�C�����P���c�Fk�����E��PX�fn ����z�����%羪��N2�$.��!�;y�p�K�%�~a��jQ�q�F�Uȣ���|E�5D�h����fj�m/y~y]&1dKS�)P�BZ^`*��?�> ���>8�FAC��<���s���������J�E�v��/��~�|��
/��Ɇ�� �ڲ//v���꣈��D����Ē���zz����)��ؖ�f�,�~�pt���mԡ�$�,1��f�G���I'�|\��ծ���`�(t�gM����A� �K1�-;��ś`�6��`���vf�l�Ҙ��ts��$O�\�t�ޏ4LfFP�7�C��Kr�(�`]h�=�=�r�07�+�����ㅚrru���ֽ��#����������&aO���t��p�)%�H��bhPzL�I;�=�j� ��<A��EEZP�;�P�]��:9"r�r����rC����qu�y�&���Z�����O�$Q��/�UV�P���N��*3-�Y	�-c]�>�\D}�9�s�k%���V�\M�mJ��qv���5^Q���7��Q��a�`���CO4������|���N�Z`k�q:4c�V��p�����ѫYx߾$L��P[��%A��Kxq�*_%a����Br��]����-������6��H��OP;퉁7d�f&T��fh�G�Y����|���F����X5���wl�&q� O2N
ܗ;���]�P�W������,l�H�|8�L�Y�8:�B���w6qŻ���l-��`)�MN}B��Ղ8RAG)����L��Q���/�R�>c�������
���)� ��=�V	VJ��sA��m������R�Mc�ߪ8�T� ��y��r5��i�L��4�X�����Ϛ0J�tjEs#�/��Z�4��~a�2=��|/���Nol���!)B7^�Ye�Fm�Ѷ��jA���迖��ú�q�)�ȅ%E�6��wc��i�D���'p�9�)�h�b&����J�k4����G�,�	̊H�f��y���Xa��v��!��/��d�1��kZ�`����;���k��5�w�B��ȼi����r�
����T��0��~��a�cK&Fk�t����X�ju��C��������D�[��c�{�9�"1\��	�/�Q[i����RQ�m�ZḾ���~[
�qU�/�4)ts���U���I6An�92�E�7ϕ�,�{���q�+�.�0�����}g�`��y�-�8Z����l2�� �}�R٢��rc*��4��l����G]%���lv$��K�f ε�M�F�����$�ܰ�W�I���t0���{�a4�=�>��5F�N-"����\1��F]�3R����-����+�⷟bz���?d�$9�6z	����6����Rl"<Mo��+���}'��W��nx�<�\kU�y��B�ޝ�nj\t�6\���n��횜W�E�P���!�B����Q�A~�ٯ��-����%��BO{3�'��2��'E�o�|�?&�!2�U|��D�(&�r���'�D��Eg"�����ɯ2\������O��O�],`1����P6WvB�oLU�
�����c�zȗ�^O�[;��;����F��q������p�M��
ΐR�M`��c�p�,c�X�"5���-FM��郙<���5�)ͭ��ұ�y��������ĚBH��_���ˡ�ԩ�-f�b�Y��m�ZM�s�e���<�.�
�U�\~n8s�rf���3b).$��0��9š������8�����>��>�b
\6��7ү�S���.v�E�O|��_(S$3��N�V���~�)ٵ�(��F��4?m��z��4�Ym#��n��V5t��Դ|���Ŀ��ă��Ƕr�����W�x�Q-e�H�C6t#n޷�6e������#�Q��m�4��zy�M��`O�[�������6b9U�������#��nv��J�����L-�=l���:[2�3�wE��ڴ��jN*��Ő�NnP�L�dQ��Î���xnDx�]0�K]$U�n��k��4;uHzJ���ϳ y�u�R���Ƶ�'��y4�������a,M�*��l`��Nb�~l�,�:�����-Jj;KX�Ҏ4yh�`/O��m��F&j��b!&I��fR���/��e� F��>�
��f�ҳڃ6e�����a��ܖ<���d7��%��{]<�D����&2�i��>O�lkм9��Yw�h�?�
1�������8p�:\�(�l�,�w�ɛ�����n��q�<�^|��q�B��[���`Ёп������4�xD��G���`e��)�Ӛ��(	�*P`�$a!I�Y�rG��Q�����P���v*[�<KT�����}��נzY����ګ�%J��r�AT4������Le{�)f-����p
Sqn��	��/yc��ur~y)ЋB����u�#>1z)~J6ݪ�0�;���'�r��q�	� Ѐ��i�$��2W�K��{˓�}�;�7��.D��ţ]S��kP��x�&V�\O��4�s�oe^+��}��/ ��,�l�xU*f ���D��t�:52�	��Wu���NG&���b���2�� ���X���5G/\C�렙��9��M�������>Z�w�����iSaw�p,��{���vQ)���ӢH��*��5Ek���F(���V�5]1�>�o9 Si�L�p��8�A�%�M�Àԫ�fC�2�ق�j��5K�[@���c��;��΍�Е��]�GH7���L�/R WĠ��ѩ!�}�fɜ��]xp��U�����q�_��/�)���c/��������|����V