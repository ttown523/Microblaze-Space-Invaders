XlxV64EB    1b98     9f0�	��r�ݠY��m����?p�N����su�ivV�^���i����z!�P���τ#D,`5q��zg)Y�|���}��
�;�����s�G-���I�H�ɱ��	qL�۳h֭6W����.i���h�A��>��u�z-M��Y���򬿓<l��B��5�	R�k��0�@0�l艋�I=U�5T�rV$�ڪ����e���p%=�i�5dS۴V�:Q8 'MaU2�Ô��Y$ �#q�c�*�[[��8�ur���F���df�<cj���񏫁`���F|2�W��;Zox���5`�^�p��4ٿk�����b���KFB�������7em�fA��r!g�c�4t3��ʂ�Z�}(sҖ��������l2�3��J�3���<4��2����"P%l-,���4=q�i3j��L�����ඐKS��f22�Y ���Z��'P����c�U�2�(��1 9P�I;�y���.�s�d||´�K,m����ܯ���Y	c8%������"�o�K�k�ϸ��������&�ֵ;�g	��~��2o&���Ď�ْZE�P�[��N|d2Fn���1��aC��פ:��6/K-�'p�L��F�6d��rxvI�z �kc��=���s�Eب�IL���{t�Zi����#M�A�e$�輾����}{�L���<̝��a.����A0��ۤ�����dEC�.����>&�^fdH�����#�ȃ�[7�MB�3��5��7�Gf�,��J�k�;�cr9��?o�hS?�3K�fbv~�v�F}`T��� �ķ��"z��+��VA���{&gG|�+il���ӻ�NoN^�rn�c�Gq��TK"d3����R�:!��$� ���5TѓΝ.�
�	`\���NS�Gİ>OS��xw������"Et�k^�k��Pd����~A= ��r��Sn$� �r�(�l��Y�1�� �wӌ���@�<���H�]�ȞٶC[�����c���rq�{+H%|�r�����Gp������c��.C��Ѭ�{�$�28�u~%\&�y���By0�:J�� �0w�]�"�'��N]�켏�{���z�%�nU�?o�]cF%/��L�\t�B��\쫷mT����e�X�!���ir�
;pWqGK�(�z�c}��#�J��Ư�������F"��(�$�lbV�I�F�6YL ��A��ӕ�L�kŎP����rˤ�*��Y�s���	�Ep��Z_Y�ǅ�=�á1�sD<�%�=���'��p��N��ᭈ�j������\ޅ��B&%[B&�9��2���NȆ|��	����d7��.Bk�rF��JJobx��R��)R?��H~�i��>z�Q"�<��=�3��|)�ǡ	�=+z��σs�d<z�,B��U�������L�Ґ�[�j���c�����s;I	 J��9[S'�jz������]\��2��Ч��w<b��'B�l�~�6�8s ����f� &2V�Q��5�}U�)0���u+C����(��n�U�G
Uv�ɀJB;�mKB�Q�	Gu[�RD�D��EE�z3t����0���֛������1��A�0�'yF���OB{:qA�����D�@9�h����b�9]H� ��u�=��z��W��j��ޒ����|$�O�^tK��l��fϬ�8׮󏽖c@~�%�J��i�L�����Pd���ƭ;���Af7�ۭ�h�R�<w��/�3�6�sƻ�Z�V��� ψu8�iԓ�m��ԜOn�Vv$����	k^вICOPn� b��ט	�	.ޔ>v 8����bJ
�1�o~����욬����`Z�\8`������-*Χ��=�L]~��k,�l:���[�MK;Z2��ʀj��1z![��Qf�BLT!|/�楅e��@� D�������36�	&fpϲK������LZ��m��5\��Ô�U|/�Cf�F����ք�s��mB�����GÖ�8��f��ӆ�I�"�ǉ�7��"��#DMn�n[�<3��;9��0��f�nVn[H;�{y~]L�[%�1��/�V,:g��c��J
�_Gc����n��>2~��b��oh^����<l�H?K�㊞"k>��5Mڸ��/F���k�	۞:�o��!�����mC�ۃ�:ď� ��@R(�7_>`m�?u��:!�HW�a0�	���rƆ��e�9����Êd��r<Nx1��e�)Rx��f�]d�t��9f\�$?��W!4|���l�|g�E���Dk�j��|AP��Y`��`������v,8�(G�Jyb�օ�z:	8o�.�O)I�Gu�^���1�$����SE( �y3�i�T}���G#�1��Cv�Q.�dy��r�
����d�˩x:�g��m?�B�E�~�~cP#�Y�.�
�(�S�����epV0�ny��N�
h��]� k\ �NC��w0�rz�AtsZ�*R3{!����$�Kڊ�{���S����