XlxV64EB    3ef8     ec0�"jwБZ>+���.��iU-&>��+�k�<��&b����
��7��eh~�����)��q�Cs�Q��B�򻰠�·`�,D�
kx����6��4�Gxet��U�>����
��/|�܋-�90;Q�=:��e�c�g �lK������hn���-;m��i*dm���#~6��#	�o�!]k3�Y�(�0�\'lDNMU��Ǖ)�H��E��c��԰��hl�+J�~ڬ;t�]J�����l���f�0���3t�#z�o�ϋ��T:!6A7�Om�-.c���F����.K{Im�f�c}~|� :z\ �K1�8@ �sQ���v�Zmm�1��7��)�%?; �O��l����+K��o�KK��̈́�%���%���"wͶ*��R�$���!���,�;���?���p`(�p��'U�;��S����X/���`eo�7�h7����l�0��8��F�?[�u�ƃ�o[�C�Ӵ��3���/�J���Mܼ۠d���.b�t�w�*��dB5��֩:��7Q4���>��u!��iqz0�^P�W�X�0�'�&'�(�����?&F�S�Mn>�D m ]���<!XHEM�2��u�[+"�I]pv��A���1���]�����^�붜r� ��/�w\����9u���9jDo�5�KZ�����h��J���V�ÿ6gy�M)WH%)��@$�e��g�y��m�.��3��;�^�I:(����d��N�W��7t6%��bQFd0�3,i�>���+��8�%&������CQ��[��h��'/�x�,w���FթZ?qYa7��H�,��v�@�p<tꇳ�䛼� GW �>�,����8��|d&y����D�$��V��2��jKI�t�_��d~�I�V�s��W�E��-��(�|f���ywJ�g�������<kά�}��۶(��u`���x�8��/���I/��%`��7�p��%߰|x�II�p*[�u�!sm��">�F�#	[Q��%��@Ii4/��*ʕ!����$da�C@�F~����仮�	�|Pof��[�FD˾Eɏ�;a��:�*��j�h.|M����;�u�-���W���*�r��e2F�"^�j���yHN�p@P�Jd�*�b����Eę�ފ�e��3![�Z����+Z�M���44.q���	��4��5ɡ�
���y<:z)�D�6ۨ��H+Ѳ��xI)��ڱ��P�������kм�6�6>�D��L(l�\Mn���8($�m���� ��{MW���E�Fg��!�#}p��#���8Vi�Yg����v�y�:�n3D����<M�a�=�7"�%�UΪ@�`��n�P7�#^�D4����|>���x���<�nM�Z��Vc�ZU���u.l\΋:al�h���Ν}-�k��X$�&Zd�+��K�_22v��ƀ$7y,�>�Z��9��U���rAo��a-ʩ�ȾԔ�ʀ���>��c�Yߚ���>5cVc>k�P%)�d�<P#,(|��z���S��Y7�����V�⏐%8G���sM��~��`�#����_p���r0��������(\rA�{&ٮ���4 ް��t%_93���6��9�sÎQ�d��p����i�^h�eLY!�lB���!f� �|ל�X�{�j&�>M�ɤٟL��n�}�S4D������IEJ��"u��/:��&Q�d�T���߿���#��%�y�)I<�R��_�o<�'RcM���(tu"Δ�g[:��ig,�ۙ�>	�^ x�=gvZЉSr�%ndC<��Y;�F
�ӈ�My�e��������_����x�wZ^d΄d��yǣ�m����[�q��_�ʸ��$@��*���Jl��A�B��Bb�����#�(p%ir����� �1����D�j�zF�<���Ќ{��k��;'bt�x,)H�ηZ�Tg��*�E�V-���<0R���/����S���Ed��J!�R�'��%Vp�J�1�A��*\|p]�x���=k�:|*uL���g�藺+�+s ��������*�X�'��mYf6�����HZ��/	� ?�ME �|6>^�B�Z*��p�<Ym�1�|&+���gB(Wp{���P�d�J��V(���lW��n�ӧ��r@G��*S)QB�s����"2�X�����'��Z3�N��"��+z���J\�#��fLw��wAN��A� �C��W����'uPY�)�
��㉦1S�Q��8Jꊁ���:�*��*$=l{�Ey<��89.Q�����8� T�2ƕ,q�rٴ��\}hfl�1u��7�X9�E��"�>G_8��T8�c�����`���fe�u��72I��WCFĺK��b3��W@�'�u$�aq��������5sϽ��*Y��?��F��~�����b�lx�Y{`~ÁU�(���D2�%�1|ǯtL�`� ��5����� ��� �xp�� ]z��#iC��n�S�s�y����\�y�v�WFΜ�TY"�d��g4��P���C��C+��k���7F(��6Rf	gܑd����r���3?�
[Mm5��W]�ڻ&}1tHv2U��Y�h�Lu�nf��5���x��Sy9<X���&u?w����) K��ؐJ�B�m�@F�?w#�̐тiiY*��'UwI0�\���`���]뻴���w�+����f�SA���[��o�+7���tBg�qGB�'A'��+�.��ܹ�N���O� l�<�ʀ��k8�sHu�/��k^�V������;���c�>�C.�v&�0Y�c�N4��2o>�(q��p�#7?��T�t6�sXj���/�-��b��Q,	���N�@�-�q_��oCG?5!L���q^;�}� �8�ϛ0�6n�Y����ʼV3�����jx4��@�~�m��UB<��R!�G7P�N�T����u�v�p�#�]�:�t֯�V��k�,L3��}[̛'A"� �j�^㭇.��3(!0Ԗ����s���W���@�����d�A>W'��"�,��F��&y!T�(��7k6B��p ;�MX�sɍ6�H>!Ny�ث�D�ٙ���U!�D�A�-���y�! �?�~����ִ?���LK4��O�֚R�9����)�I@A�&��(��"s�t�����Y��v�����v�l��;Ur�V��Ԡ�A�9�����R	�����o�b�,���&�G�ЄFÄ���xB��
�y�7n�� ;#C4�٦�.�u�f��Q�G���%����ey�LQd�z��a�"&�l�.�U��p�ǾUJ͏�|*�0�J� ДB�����N��0i򜹔:�cH�)�����e]̭ft��	xބ�ę� �Ig�qE�c��=ՠ�,�tv1���J�h�39���0�\���$�5�W�싯m��nkha¸�y�w7��K#�@�:�����bq����L�k��U4���^��!b�j�8u��W�V�j�V�	po��2���
��3`W�ȯ��*%����A�upߣX6ݕ},����H�hg�]�3KSVG+���%�3ǃ�����F��'	�hrs�QU��^t��Bo�'ouD�T�:nt��8ɣf�]�"ׂ�38�bG��S/����p-%�/��c�0��mR���vؼ3���P(��-�i����q�Y