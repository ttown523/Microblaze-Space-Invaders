XlxV64EB    4a13    1100:ͪ���㪕��qpl��}c�J�B�׆D(�0��^��u5���y+	��~�dX�����R ^�96���A��Wâ`���FA��`k �)*ҍ�]En�p]��( ��lz3m]$���Yi:�Ȁfxo���Wb��y�,
Ț��F��#�9��4>�_�u��T�r�X`�k�V�pj� ��o�z���\>(}�-�&>a1�ў;9Zr�q"V�wYY\����l�c�D��
��w�7���E둱*�\E%`��y����zvڰP�X��%�jt���#���M �\0 s.L���9.�4��y�Y���X$�`�۷����,�������L<���-������	���5�1K#q�t(4��K�h��O93�P���zJ�4(��6��u|n��H�����Ps� ���)�^��yqn{�~�Q<��F��M���@�@1�Ƚ.�I/s`�y�j���D�TL�����ER�Ε�.ݑ�J`���䤫Cb�2u�&��xA?���S�����cZ]�zY�O��� �0I��]��M��#-�� ���%�~�״c|b�X1\N��w�p㏪y㨱`+9ݕ��*
�dX��}��G��<��K������$f!��i;6|*�`H�?kD�OW42��2�dksBs�=qq��>����h�1CY���a�0�
�We�-M͌O!~`��FZa���A���5=-m�:$+��>�i�������4�V0�eo_����p��846�a���)E4���E��-�5
F�÷�c�IP��ĖJj��'�gfN�u��tS�$<t�xz�-�V���1��*(�v�������z43���pex��r#M��Q(�4ي	`�p/t�A���mBf��B��tn�<�C`�P�U|b
��~�6�g3��Mm�RUF�4ideմ��
3Yh�y!%�`yd}U��.(��n13�`���w�j�;ci<���t�{X�Ͽ�2��<A]P<;��[�-:�U��|���-U�]���F( ��IP���B�����Ȑ�[�LǠra_u�Rz�(��뉱Қv��M.��%!n���x��q��^�]B�a��
�R�E4#�
$��tl�	�v9�GP��
�d�h,�-�R��%66�1`^
8�o����$����K?E��k�>��;Nջ`{dl~��n���4���s`�^2Yhx�=��GԎ��7�w;ׇ�젃oyG)x��w��e����į_X_��5�b�����r2�`���v�_���2Fs ) �:���K0/� ���{���.��l��A��m��&N<�]Z	^b�
��yÄ8����½Q���q�ܯʫd�e����Bp(�E^%#*U�-pQ��`��/�L�B�s�/�c��;l԰��-X���?�@�-��(���
R���M)w֔n��ό�	-0�ABbߨ��ufp��b���6�&5�'�*�na.��NO�m�Po��;�e��J�� �_��<)d�X��7�M�|ሎzj^L���{��dZԿ@0&����K���1�����v�bp#O�l>��� ��f�$��+�|�=s�@H����=�d-9��,�Gb�?C�V\����Sĺ��u�nb�����b]�Q�X<��HR=�Kƚ�2x�o���Uб��Ԉag�?sݭ�GX8G�⍭$&l�vf�YS~�m	a<�7���U�"1��A��ޛWcڄf��Y��w��z9�լ(�,��qA���Au�#����4m��@���r���lϚ��:�hL��೨ �v�;��O���ۄ�������ߡ��߅���p�J!��p��q5��σ��"1,�wJfC\ _��PUJd��R\�����o�
��=0P���B�|���iE���"Jg䪹n�����s�z��	�~KI�?�v��x�ӹ^Ι��
$_M�)�bz��~�_jޓq�hL�1+_~7�OAIs���|J����o�4*���c�W��%c+m~c����_���i)~`��D�)����M����N�CgG��Y��G��5w�������G��uz" ���!Vw`{�����{��L��u���kM����ϴ���;��ْ},��3>YէC�#p_K��&:��������`�iI��Ũ\��n�� Wj2BU�<6����%���9�i!����>5Xpq)?.�~�ab��=��4�G�3�+ʥSU�IL���'j����@�!Φ�E�(��Δ`���}K�,2�G���&�|󟶢�"?(���^����mbt�<�7�����#U�*ڗ.JK�T@���K��=�ܦ����db������B���VtG���m�^�����Rl�|��,p���	q�E!�*�[��h0G��^嶪���D����2�*,�9!�@��z�"�������|��gĀ�څ_��L,��ms��mX��4�� w�v�ݴYj:~?I(��+�B�7q��Д1��.����:��Yō�.�7o�ީ��.I?i�����g�5�b ��Q|8c\J��爤O8�T�C�|F(g���P�i������%��������h�γ�Q�3�z3J&�����k��c*��)�#�Q#��-�As�n� ��~��b�u����t�2p,sX� ;3�/A�/���m�㌐tu[!�?�Sx����$��65~b�-).]������0h�S��ۢ��-j��F��P$��xq�"��M� � Vԉ�д���27��:U��&rZAo�wT[)L�1� ����л�l���PDK�7���ss��=8X�Wat�t��4�"�J��0QD|z����i��/������;�]t���c��B�Hj}���<1�ݻ� I�`\���v��%F�a�~�w��-h��yLҵ���@�|k`E��
�������ˮ�J���%�VbL��[cZHV(��R�������?KF��k�֚����E�Q�|�K��9��F���t��M��[���|�����-���2K�q��׀� H\�jܪ��RX4Ѿ2�xw��X?K$ ���r� ����cAv	�x8�/p�+������d�X�BPe��q4�^H�e���ʋgF�_܅��EReh�kg��W��������'9���}��rS����2�l8��N0q1�M��+[�X`�#�X�;woX���Z�ވن[��Ơo��U�m�z�ې�t�"&�YY�ESZv>n�!�z早=����f���<�w��1���Ė�~T%��A!W��BP~Ǝm�(����P�W��n�R];`S����$�P�8�V���)61��N� ���N�|��v��Q��+O9�h����ҹQCG����D;B:Kx�,ukK�;�9d�l�[��Ͼ��Kz �*K%�QX�6*���c�f��dc��������L��>�}_���l�>g}��uwx�Z^���vZV��e�Zp5�N�b�OtzB
L���z��/�/v�?*&frh�}`� ���螺K��L�������[O���-;&x_ՆH�q��B�' .�[�V!q�PXHbV��y�f�:��ۖ��~�դ���$����Y�D<q� �����L�o��wZ(穄:���/ywj߽�6!�JF5�ڙ��4s9ۙeC+4>~��{h,�@���J��ا2���G��_/h�ƞ�p;��S���IjKE���aMq�Wv�.c�&{@\�����iz��|���0�D�Q���(y�z�l3:��R:ɰ�����J��
њ�����dK��?��m^923h-pk�ԕ�%��Njg�j�����!EE��'�4���88�NY�CX�~�s���ڸ�ʥ��D:
	g{�_;��I",��y,�BO�K�Õ�*/��@}�,��C5��N����� *MD�[�!��>���yД?P�8Y �b�@��7r�z�?��2��W7�;�>tk�:d�~or�7>7�Prg�#
�I�l >u�N�m�F4�}� �����Z ur��(zjW����������9_�� ^B?�9�A	Y��e=ʯ��Ȑ��4�8�)���U�1�؛�k/�	`���;��$��9� ���`q��Hʞg�~��lK�
W�f�_����.�k�H-��b���"�����Ѡj��R��-jt`[T_eP�^T;M�SI*z�x����L���1��QtAfsN��L�et�Y����1�
�7�W���e��|:��+�y�t��	�<>�4���Md@ML۽*�h���1C[��.�$:���5