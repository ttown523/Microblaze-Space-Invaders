XlxV64EB    43b7    10d0� w���Ρ6:\�뤥k��J�4�����v˜��6-&��t pI�r�)m�H����N	��� f��)���$��k��T��t��~�r��7�ᰆ_�.ƗN9�x1j�,\m�#
Vt�Ω�D��SC���Z���H�T?4L��0�BJ��]����7�S)@�lrgC|n�N����M��Lcd4Z6�������f��	!�8�L/� �ʵ{�� ���э4Z�|ב	N�l�1 ���͖������b�&��푼�	"$f[������[���v�_��yv�1��hҟ�y2�;1�R)���%�}�-�L�9�cϚt@p�YV�V��Xx�_�O��MVwV0���W��2���{(=�kAx������ާ���u�j��`�Y��N{�c�IS��T�i��vY9o�uA���᭨,�H�姫}l�jZ�(ȕ��8�@�I�_�<����e�䘐�X7�pa�F����@�3[���v�l��p�XĮ!���O}㉗\����`Z5��ak�+n�]�zg�x�`x��Ә\�x���G�[�d�)z�GvZ=����1�����?A)�)/���+[�j0�
�A�m�dX
�yӑ2����ݽ�{W�* 1���c/�ŭ���p�m+c�[V��6�BI�2�jy���O҉�%68q�I��S�$�)�y�^�mƤ��� ����������n���n� ���	o-���k���+���<�mx�³5>���lN�!�!��#��Dzᢪ�8�3���p�� ����e��{��y��W�|Ugƹ#�W���* 3�!z�m�VK3�!����鄦*�u��9����v,M�
N��a�	,A��7测�g�Ϥ��S ���q��з�
�XD{��AM�$�v3a�r�J:���ql�41��ǒ��/���d���OL0�i�N�@i�9A�����O��ιVg6�cq����1���״
!�����,��I<�]���m,ZB�x��.E�0��UT�n�nF]��rSv�,��Z*a^Q��abbz���y��[S��B�y�7mi��Q���:t�S���!B��:�QT��D2&e~p.�pw��=����h�a�����6|��G���[@D��8�o��u@/H)�%���V;b�c#��O�}���}ҫՑw_�Y�4����)_�C:W([.�Ҟ!��[���Puv
�� �ͻQS�hO
����WHy�)�|vVsF~�c^��U�F�(��[7�U���UO��X)���B]�,�@U*�m2
�J�_fB����TP#��?���KI4�D����?�༑��*8k�f6Y�t��:R���g��(ӷ�YbqN^��V��]~�C�"O�'f3��-�C�|:����7m17.bc)r�%Dק*�Z��OP�1T�e��_�_�KvR!� �^��\B�<�:N��H��䄋������,�D]ג�D���Dܦ�+�!"���+��q��Q&$L+���l�T�ůb(���ٲ��p��Q���&�f7+�������&ĎD����wv����g�� ��?�PKAk*���T�ۋ���S�����ǋN]�\�̏�T�9��c��	�[���v�ӗ��w:$����T�ˋ�$rj�$(T�2����6F���ut�q`A�8pw40R�"�	�ע����O�����T��=9u�  sV�eE/x؆�W���W��4�T��pg�O�o��|Czn���<MwV=;_Q��	0�.�d��9h��%��uݥ=��� ��KYu*����ϲ�v�č��LTl��K�S��+t���r�S��r^�]ms>�*��+�wG�W`}�0��
�C����Jړ�2�7Q�Sm��f�>�/��_���]�����>�*�=������&�6�q���=�ӂ�{�[/Ne�5h|��Z������
�Y(i���0B��=�J�}n��Xd��[��LQ��cN�L44����
V�%7y�x�
=`�Jv��T�Ѧ�Yo5�{lg�v�a�l�x��Μ��?T�/!���`Ҷ]ޖ%�4��W�|c�/b�˲.0�Q�_#m�@�R�Њ��~uչ�dOk.b�r��֗����v�>��F��D1�H��cC���i�Ñ��@0ï`��f�Ot���W�K!l��X��N��=�<݌!�E���a�>P���^D�����zEȷ����R�
u�f���]/�� '����~L3�k9w[-�����"6 �a��W�=�Ah�!�Y��@7��X����5���qf�w�d߂��r\ }������A
���@g^��.����,�x������Fq�C��&�9(����;�2�r�TE�ca�VB�eT��0�������p|�|�� N�r?7xk�\�)��"����(��$�u��[+��p�("L�q�TIqJVR(<K��{�5��2�r֑�&E2I�1*�Q�L��Z�>�vM�|XB/u)��*�i�T���{`��*�����	9ј���m��>EB�枯�C��s^�頋>(AC�a�c(j��:PQ� #�y���@���LK[���D���1�ٱ���3���%O�&p��5 -e}�0��`
.bA�vȈZ���e��t�O"��(M�D��9\�K[�8	�c�H9���vJO����<�8f0Vl�DC"��l�s�Sww3@U]Gq^��mq����Y�n�oZ���ЈF�\���bxk���c�w�ٰ*!	�U�" u�4d��P� �e�W�q����U��0�k�ol�e�"{(�q�*��LV��y��i�6�!�-�{�a�ѯge�ٮ�1�ol��fk�Q����T	M甁U\-���M���b�������\��^`�������{l�[V�U�}��
Ɓ�(�4IO���j�t��>b��m'���f�Rℯ��&�
`�����E��FGd���	�b{S�{�r�����ۡ0睍|L�[R�v�Kj0����,��X3�˗�=��g�`l��e�Tu1ǓZ��}_e�o�IA
�D�����ܥ I,��P;�������FQ�c�!~����p/3rEu��9����6�Ji����B��M�x�Y�]�U^�.W���qe-M�:�W94�o$
up��s���pT<��E�M��&Q��?c��]U��AȺ����\.�t�7ڭ��hԓ��z؃��'O�!�~5I:�qAQ7� ��)��έ�Q%R�*D���"=������7��V�E���!��+��j�����d|�,���	q�!R/#�(V	���ZB?���@գ��6�vB�(�"���=���ަ����e��ޱ[���Z�M�,T�S�"����|-,�n�A��f�o�`�^W?BY��Í_[�����O-@�Oט!�����-66��v$.*���љ�|L�)m��:���8�Ĵ�X9&�쭯�� K��f���Z5�wRH��
ܻ9��F����:` �?�o�5�#�����`ӵ�d66W�U��* }=��Z���n�~��S���Ȭ��WVF��વ��O$�H��Zf�%�#:�F���� �1<���&��b�.5dS��`r���������f�|��L����a�C���i0m�y�?rYa���MN�>���V�ɫR��c��G�
���#��p���l��vr�I�\P�+K�����?g��jww�7^��;H�/��ٛ��N��h��(��vZ��5{~C���a�l����y��b{���C�u�}�[��lz4j`���d���I@ $G T[?�߰2���xү�U��ȏ� ��v3�Q��S?��P���8� �b�n������)�p�D�3���}31	�1���~��Su�i���6�T1��jwgj��T�TL�P6�["��9��wA+�1}�Csu	��Ne��bx�9U�{K�ж?̀���S\�߰���0�!t'y�6|sS�1���뽊����4��2�+��6�Y�R��fS@��`Ӛ��˟X��9_��9�]���Z�ߟ���omw��r����\ p _�q�D��x����b�K}F�AR���ϻ�:�*�ಭt|?{�rP���L9�y�Xp�^�.��KH�`���1:��h�g���2|�Zϕ�/>�y����!b�-��q�u7z&9�L�t(��W��ỵ��>�E�Ep�+7qVw��ɕj�o�