XlxV64EB    2232     ae0����$h�9�u��/����s:���->�/�7*�}�"Ryw{��~H9�ii"�?��$XF�38�X�A�2�e��V�Ra��!�m(�/|^C�w�[1���6�2���ѫpv��M��� ��_�n�˄z�>�V�1n�R�i~r�u��}�I7Pv���cN@�Kp�Wb�ۊ��$^�Y�![(3Y���,�S��ӜhX�S���_s)�(�6����-�R--���	om^��*l9�a*e�k|�#ȏ�����e������cP�����jڗ_��q�F�#��\���si�T\�4'��)@{��`vuf"W�T9��8ox+��>a��_e��<�A���[~��ɇ�Һ9��9*1�M�_��_5�����R��+���#BE��8�	� $�w���b��c�a��B^6c�]�^�T�v������TkRSb|���{����?<`V��n��/ҳ��:����}����6fę|bZ�y�̢�òO���vm����ؘz�I�� ���D�҉�λ��~)�ܕ�Ϭz=�Qճ\{�ۄ�@U&�G�{%匡4�gb懨����!M�!�\I/o��q�S���#4�M�Yv�1�فK�hv�d��;NK�9S��R���f���r�@Ǜ-r�>�x7r�lv���?�ٻPm�h��m9�5d���+Ylي�mB�O��ŀʪ�a�ov�*
L؅xg;�>[�{1��4q�R�<�!~�2�8��������>���b!�v�-��*�����6��)��;N�	$x�edFS��p�� ��쁓��ZOUӅ+�����dX�m�5
w;}0U69&��������e�_	�����
�X�>�Y/��	Z�h�e�U5�fц�M�MD���� �	?�y�l9�BC��e�����tI=��W�-�>J}��ȃ~�6�z��d��_��h\U9b�8�����P3G�w��1�V���(��!9�һ֎Õ�b��Cw˔�	}@	
"BK���c��)��S-�g#�W��� }���iN�s�蠔-
�r����x��b�XP���HS�0��5����a8e�d�wuu�� �i��^>eB��}��Pڐ:���B0rʝ�wݻ7B|�W�T*��T�Fc�=X�^�P���S����
�_����|=D<��;}�*A�'Z��q�1���czG�L9IҴ<ƺ��:U�ɳg(�y5���〺�\����Q/�u?%h,m�����|9��K�L�<v�$�`�M,]S p����2��,)Y��,q����ԁ��;~VkǺH������_P�YA* ��L�Ց������'=eK̀#F��,�s:]x�0,(�5Ӫu`�J\QOᔼs>��e�''�����`�&�:�^��'K��q��N����C�9���,&��B[���i�~
귒��ҾRX���wX9�o�����Mb�Q�|�O�4?gP� �-F��a�:Bp�uu��l(�fW�2�����r��i�F���h��_��@<τ,L��W�o
�U4�����{OmX]�9
�y@\�}�m3L���^~zP��KJ^�z���w��%�p6eD�K��|	�Z��R�:��s��ڈ/2�6j�^��rzΫm��1�>�)F�fWQG�ү��p׾��u�j�̦���ؒm>���ۦ����?"�ͨ�8?��;Erf��`�C��d.�D�5e���PsH1.j�>��uG'h��4��ޛ��d�ͩ
���9�t��C�lx��*t���i-l)��=��Wqgk�X�<f�%�JC�MI�� ���
�G�i�]{E��	��}]Xʍ%c~?���?����a�2�~��.��ɒ����4��Wr�8���e�\1� ����'�/�|���=@-ͯ%`��� �.Q@��jm^  ��ۉ\ r�x$��$n,��I�DJl�Z^9y� ����[ܨ_�E�ΐv��C�ٞ�V����p��g��U[%�p�=j�{ת}4Gƍ��m��� `Wc��f@�Pv�����LF������o)�* �</- h��f��L  Lr˿L���Z�v�ـ�e����W)�����%���k]��"�o����2�+��>6��`�N�P��."�E�s��Y!�����$^!%EmW���e�W�ǿ���9#OX�8��_�{�fd_^�`��������x�&�QT�,���I��Q�r�����^cߥR��� �&�����G	j�5�甖�W3�9P+W=����}�bΪ�5�Ƙ���U"E��Mg���D��|fK�1���q�'֮�C�դ�GrADY�?��3��ɕ�wU�<���EE_-Ω�$�-0����*(ȶD��U�MS��!��k�T@1�H��Á%0����V�/��W�1˂��440���Ә�;�Z#���vX���]�X-:��2�a4ۊ���_���6�?5�]����-ɜ�u2�0��}����/�'=*y��&aX�9Rk{Ο囱y`L0z��g�kZ; ���02r�%�TҨ��Gn��y��K�9���V��hX`p�T�jE3^ښ)T���4�++܊I�*rbўݤ��ɤgx��%s�+���*����hlNz_�}$?A|��yKN����طDW�-�7Y��r����L�6�� �$eϖ����Y�v̈7��|���&���;�ޏnEAWT{�}��|�U���GV�Ox����))c�@IՐk������O�
�BR�c��Ŧ`�J�