XlxV64EB    1648     880x���]-@M+*̔[�r�5<q�q�I}�p����C*�G�.EGw�o^ݟ����_����n۹1!J���w_k\~���BN|N������V7]�b���6�C�z��3t���Z �M���q�u�ж��P�"xC
@��vf<�d�#{��K����*$ME���"]Od&��2u��fQ����j��xNs�O	���˃4<�ޔ]/�rh�Iy�f�o�Ϝ��k��#R�w��-c�~�]��nP<���tt�ý?��Lb����ue��p����F� �4�9��y+������q �^x���+����V��b5	�Я�e���Q�U?��-����r; ��1����7N� }�ݝ 8��֍�a�@f�$1�:-�Qˣo��u��{J�� ��H���"���AimU�-�o3����C����+L󙚄�������JZw��G�{(��$�0C�|��I�J�y��$C���C���ߥ��)��ܵ[�%d�:6�jH�&��ia�hh}�U�V�֎yi�>��I�e1�Yt�)��ct:6OF��@Y;Z�~՜��.�MC���WQ�A��D�]�~U+g*���	��MI�?X����P���g��Ƴ6C7�"���R����c�aT��BUB�pBa^�<�{'���@*�<�/k<�����2@�A��� 3�C�rڲ ;�l��zQ�@OaUTնC��,�G`���kGeOb����~��<�]����v��Z3�Zm��lӓ~:�èT���:b��k��4���:�۴86^�a�7���+�5���D�7~���m7���bT����{�~���J�5�n=�ފ�>�b��K��ڔ���g�	���~9�ٱ���Pѭ�y�jUˎw��t���|�:G�zb1��*/��ߪ��A�p�.W-��x�F6�J�l��o���W����ɡu�Rى�����w���s��9�	��Q($�G��W�-�󎨏�/W�QT�z���!T4�lGm_�������<p�o�d�J���ȲH
X�҇��r�m�lN�)Wӵ�$(/����"�&Z���x�7��~�Q�%���8Y�����IMV7A-��2���1<Z5A>��V8�
�d�n��&r�.�=��:�m�h6��ح�p[S�Z��-	��+qk�$�"���f�%�˷�y�ƞ!]Pc(z��k)r�H~]�_�)�$��X����
4�\"?%|A�a�aƾ��f8ŉ���rP]�^���MY'VU�=S��%6���������Z���o>t�X�{��t�܄c�P+x3�R��������2��w0��@�&��<�7�e~�k|��g�ګÝ�q�-ý#>�u|��Rk�N�t��������_��cL�O��k��W�B&"��t�B��RQ/�/�
܋����!��~��{I������z|G��m�՘h5�SO�ϰ 4�:��Jg6�[n������(2����[�@��|��ڧ� �\��zςt���[���8�6�ۮ�Ƌ
zv�~���/W���.�+ǹ�?=�͜�T]
�춌� a��X沵�w�G�CL�60�s��U��m��F���Y����#ٗ�e�c{j./�)������a�����5��@��0O��uȏ��GcrCD�|�;���l�r��I� z�C(J�Թs9Q��W�@�Z��%�B:J �@4̓Y	؊�ȯ���k�f��^d��>34uB˳e��ZC��,���5�F;��gݫ>�OJ� � 7��S�}♂�P�t{P �V
����?�އOeOh )����T4�1 �:<���N3�/�۫�4��AA.�z���,�-������ө<z�u!)�.��u%O��=��Ҿ!�P���{0Jb�m����]|����C �� /ِa��K�ԒonNL�����l�6y4XуZA`��V�㸬�cƯ�R�L$j����u�Ju�Ev�����9L�~XA�JS����f�|�a�Z�N�允dUL.�PR��Zy0d�b�������	"���3�}3�s���ʎ�4�лFP����-�
�K�4�Ꜽ(��ea�T��?�j���v��<�?2	������o6�}�h2]yd�!�i7吟M/ �Z����B