XlxV64EB    17e7     9b0���&QA��y9{F�0��E��C����*j���U�9�����D���]���؂��;uQ�����Un��}HߌF��~��۾�lC���q��(������ߕX+ɵs�bDO�����	/�71����d�g��^N4wp�Sl]�D�屚�m��`R�=�-É2_2}qWМ��2�����r�m�EH�P%ox�>�^,���4R�ܾ�FR8Q�^{?&��[UDe�x4xMo(����W��Co�;��[@�V�#d�1l�7�+���6E���|�/ta��U�
���Q.�����P{�VWV?�ͬ���)ZM���d{��3'U�
�Y�)f�ָ+Gy{�����5��}�WIlU�ԓ��ݜ�d:��]��j'��cW�:���x�VM�?ہ�� �n��=:{�|3h�juN]�I~��{-��_ⱊ q~\��5��v��d,`�~�^�S��n�W ��7�EC�ygܶ$n�>��1����C+63���9��JE���mWq�b��ί��?
�,R��<�A	At��H�s�r�ƁƊT�e�����_����<�[�ʯ�M7�^M�ֶ�%=37�`y��ǰ&]'�S����������T� al`33MV�F�M,tɻ���m�W����ڂ�_�b1j�,�{�@	��rG�U�u�V�]6�ҷ�_#�,�VL�7$�r9J8�����ް��dSb��d�C��V����[~q�OwH����F{�|����^<��(�iF���*�.�=���3Z*��A�uT�N'�e s? �\Ex�o��f���'l��]3��y��u}�`Q�l1I/�/�@�?�՘�	O�pe��ѵU��r��]�)�������{���7�M,�J�U�;�2�!T���֍YK'+��(R����,�%h	k6��q�s�"N�54-�����S��^�2d�]�7 �ǂ\7p�ɇ+s-[�,�m��`ku������Lt�K�.K���#f=b
}���"�1�l�;m�/�
�����pc�ɟq����;k��D��~`���%C�h3�¢I.jl6�A6��g�Aw)�4Dc��]G?|�>�Q{l* bj����D�iQ~�{d��U2���=���
	�����a�a ������!�8!ߔZ��1�R[��`{��n�Μ�S�%|���#�B&\�<:h�y7��u�
X�e�~��i;�|s)^gd۸2fj��a1#�R7���B8�(yz]���]�O@j��U pK��bF&����a�o�rs�f.[�������'�"���/�כ��e�Y��g�T�r��}lɤo,�����ŗkDF��<+\�_h���M[s#��f
��+l�S��X~�K��b���>zK���Yǁ��>*7._�҄ �C�v�q���"�{31	���m��,43��YX�`{�@���Mx����O��\s�e߆���4M9�������0���TL�;��s��,�n�v�^�G�9Bo;��@��Z���n�A��JD ��O�D��̈4���5�X�4��Ze�Ь�gNBh�����9�u�j��$u�r��pAXn%CNɼ>�.��J_ҏҼ�kf�`�$s-���K^��y�k _�ǆ��`@o�aý�E����ۯRO.D�����gVu��J�d��a�®I�Tt}������y���:H$N�+N`4K�GT��ď[���(��m��dl1-ͫ=���1D�)G�D.=Dd1���
@p�l�H�TO�B]gQqj�wG�id�-�AՄe�R��;�%��:I���f�죻f	p�4��&���d	Ĭ�~v�����r-�s9�+4�, ��/�y�!jՎ�����y��⍙����ۛ���%��{(T���Ga���j��|�M�f��1����w�Y��<>a1E��B�N�_�4�R�yNϴ�CYC���͗�k_H�,���!�w��7�s�$~/����ADTid��C$����־JL�;�m���9�x̑�j +���ύ9M��$#92l�#���1���]�1��=������˺ޑb�����P�)��ǝ?�	��WZ��
�w�K���-ղ�\��j��}g�
���Nt��:�A�(�J3��h9�L���AT���n��� ���X�����2m����#���wK�+{��l��#У�%-�Ҭ
���� ɮZR��|��M�Y�`ڞ���szU����l���p�8�L�*T�jm�5�U�� �7c�>"@���E˩���vV�jt�>�ӵ�??A\�L#�e>���e�e��"FY> �P�gO�	���rr\Vx<rIa-*�8=@\<v<��s��#3:�����K�������7yAi,�
�rQ1\;W�6^������wr�/9�5���r(��_㚺�V[�4��<�