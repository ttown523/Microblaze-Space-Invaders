XlxV64EB    25ee     bd0!�!<=��f��S��(�d�A�b�vc����I'������$�)�5�YtP�Oŷ���֘ ��a^���K0��<�M	���'G��(XXFe���,�� �X�9u�a�gAc}Xjy��eJ����;	8�=��R�fy�n���A�GpE�`E��*�ڴ�t���Bk��đ�<�(��K��O�b����ގw$�3�:[-E~W�d���0W��������LI<��@4�I:5m��|BX3\f�ލ����+S��m����Zz�`e9��^��yу�3�+�9Wdo�*o;U���)Xh��ܝ�5`���ZԸ�	������HJ������?�Ew�u�;j�_�0N��7e�X
;!k� �߉#	��@#�Z��p6�O��<=�i�Z�?W7+6���C<F�Iy@�����,��h�b�]��5�], �]b/kO�ѲRm�G��_@Ʀ�8��ͱ�c�H~(镶I\�
ňU����Ȯ���3ځ�n|�8i�*]?n1�&��^1����z@��Hμ��qXӬx��>Җ�e��R��
�⻇�J�8[
�#�L��	�8�*�Ȅ��Ƣ3��Bs$#�QnX�z�;�v�)�;�.�u��~]�d��_�d��O�!js���p��<I�6&W_�<}HT2t���W{_R�!zd�M���%���� \լIv?��f�3���gj��c��w�x��,���\�uy3 ��c�)l�J����gZ�P�1�sF2l�M�y�n"�Azk�*��*�<])k�������#����r�ǀ�ؼ���eA)t,t�u7jJ��A<� ��	F4�:*eC�/��*V�М�j�$��Dq�M�ؔZ�@6�=�Ť�Qx�$š������J�ݒRAvѤQn<�y|">2�fo���:��g=[d �K�H�[��3����Ȳ��F-S���Y�f��ɿ�y�)/ڀ^7�:�φ���8����݄�ǚ=
���-�����u�\+����}�J������}�U�*w�4X�\G�bNY�|��)�6;�l�_�DM3� �#�2޿î;Q�%7I6�������Ed�@ZwˊnE(Zz!��[�NM�Ӛ���`��]f���Tп��k���&����7d{F����ԝv�V�V�G�M�3<-���v#vnG�0R��#�X:��ߚq�^,����{�<i���)�6����4W��y���#⇡H�~�:<}E��0^*��@�V�Ùl6��G��{�Mr�ȅ��(���h���3�jT�e����(��4[Y��CD�R�9�T[�6�E�A��F3�,m���6���Ɵ.�����T��vs�y̏�e�$����H6��� 1k�<	O��>���<��v#vd����.@�?�w��f��s�~>��ˬV����!��x?�ص4	���B��B�g�gX�:��{Q�� �l�<R���=��|����k~
]
|řa�9�T����U��7,@���G�ҹ����נ�������:|���Mm'���g���
Uݖ��G���BF��bu��?ӡ�99o�_S�����)�<��$�Ȯ9�`�P��M���n��޴z�v�r��%�6hP*����w����흯(���;v���)T��g�/�G�$Pp��s�m���f�I~#�p� v�����1�Tv[���-���jd��k���`��	<=��1��8_��M���};���t����1�5z��z�cq�%�~��I��_//�;��T�����]eN~�)]>�M3�x�[�m�Ќ�ӆJ)�濊u��
����9U]����W��Y?�^�a�����U���v�����=]�#���fٱ�+߁�8�&���R�Jf��ɬq�׆�uÊ1�To������Vo>�j6Yfk�ȡ�J�n�\"1�����S�aD4y�Tb��y$:�E�k�v[9���,�KΟՙԫko��j���L��u�LEX�����#�7b��$���9�W^^�*Cy��Iqf�8�y��-��O�R�s��
��J®g>p\���Wu�I���Q�a��F�"mg}R��1�x��>U06p �Ӫ��B�����~v�o`Tp�.����rk!���Ж8b���ܚ
w���a�= �e�8EqH^ED���A@�z|�斬�-�D`O�N�&��2�{�-�0�X%u\��fZtVi$��ׁ�dS�(վ4�@)4��6��2�l^��0�"{��GAh� �5���M�ߖ�é]s���i�-�N5ܧ�S��gu�	���m? ���\�����-|�Xr_���Cݧ[�O�ߤ���Ǳ9#�M׎`dhE0�����ũ{^º:�<�s�c'��1]7{�џ� .!=��0��͡�Y	g���b24��VQ�J��5E�P�B̊��|���>�V�w@uTF�~{�5�ٯR�-����tx��c�B�a�l�p�2X��(�@���fR�ԡZ�[�x�C��*f�����ќ�Q�,��VC§@�>����È�H����gˤ�����*N&���b/e�ݻ70���T� ��Gޙ�[�lH��9Z���i���.��D�0Q'L?��{��J5\L��=����.В>Wg�y��;2����Y���F�t�6CںY}������z���F���F���[|�]�+1����ɯ���aq�'�e|�!�d�5� ��u�A�i
���/ߕ` ���:y��K�*�c.�)H�~��� �P����ě�7�Y��b��iy�L�Ӑ#��sk!'G'0���J�S���:VUj=�m�
�<�>�-Цz������1�v7�e0��[���#c��Ϫ�W=��EZ����Z�IE�����͂P7h��zU�x�h�g�]�K�Ɵ���&s/�������������mA"'�+	c)��Z�z:��rH�g]�����i)4����v��e�k� �