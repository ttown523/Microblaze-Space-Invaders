XlxV64EB    71a6    16f0�+9���!g��r_���xQ\6fY�w���{��C��)^֮�>TLe R�!s�.����W�( 	FD����yy�W�2��~�ܳ��)���X�#2eBlͰ�o�Ag_f-&�yq}Q��5wNTC��z��J����*����H(�o���p�p�H�'����8o�ъr�Y�_�,�?kov�,t=�)�3�"�&�m�2������Cy n��/� �L>Z��.�ʙ%* 6�M.��/V��k4�9�l����a}.YV~F4��"d��
��XD<����%��'�K)����1�>Z�u���j��Lʀ��ϋ��湏#6d#���n�
��>2��y4Ym`�#v�7Ժ�{�c�X[��z��-B���`+�5��������<^���ǡ�R�?��jf��?3k��P��/g؍�2�΃��g"^-ے��������ni*~��������pYk���V�-O��6��Y�l�Y�5F��8"�Gbzvx������;~��֣��@�
ޯA�r��9�O$�;�<�+��y#V�}/q][�3���:�,���Z�>�c�M�p1�Nƅ�o9�%�O5�a���Ap����oF]E�W0�R
HB�WR�c=�����	>�qR�֓��3N��T�ƽ-_�'�`�3��?�*�i|����,���/w�|��n'�c;��Ӳ� ���	�:!t�[��@��9{����=�ٶ:�ro.�u:�k������\��CD#3�Y��>8���^E*ʦeƊ@7��d�ȡ���=~�C�ڂ~c�(�E��|̕'�h�����]8S챹��~�,�Q.�Y-�z-�?$Ք�e+�T�T��9OU�eVDI\\^�}\,Q�SH�fK�>�׉G?.U%��o�?��2?�)��E�j�4�iH��{)��If�X�8���v_e�,��/��p��ԍ;gߢ�n�3����,�n�lO[�yM:�*�3eXT�$�o@/3����ڸԑê?������YT52a������Q.;��І�����0�"�����R�;��bl������b0)��P��)s��as�"��O"<�h>ö�O���)U*|�2sü��aCX"�'�X�uG��*����ց�a����E^�!&ۊ���).����w_,�����7�-T��ֿwΜ�B�6�;���F��ND!���,&N����i�o��Y3l��ʿ��iٽl�@��
Q�~�{�t)�Q��A변�q�߫a��6�6O5\��[�W�-��*�0�+�ڻat"�ΔN���2ˊ_=^R���yz���f�O,]�!���R�qi��ʽM�)�v|:C�2����_�T�R%���0_oh@C9\W��a>ES:~��;�ǒ�_�����fJ�^����
E��r��zY!"ǘ�s�����vB�h�H�婐f�	�F^,�VSXJy��qOǮ�F�#�ǥ#G����o˓��-7�e�ӯe����/�� o����V&1$�y��BDJ+IHt���
pƂì���V��$����֌n�M�"ô��j�� �Zp�����4,�WLZ���fM���ŏ+���̹z�d�������q@�9z`0u�1�%�)r�:s�#���=�=]�����
հL�$C���l�t���2cX����/H���VNm�@�u�!��E�P�h��Ͱ��M�҇�W�S����
�B�����~�^[�Z�z]-kx�^g.w�˰>F�Y�7}��Ck5c��4
0��c�}���Y��zːU�~��n<�+�f����w���;�YST E�TKˍ���=���|T��es�<[zz�����"끽à��]�wy$E�P������U���O��*.�Z6C�g�9�7��Oٱ��'""K�*b��&]��V?�a�I�ͼDb��_�-I^�8OAl���xQ���,�\��'�$�͘KG��i�I�;��8e^��;�L*��z��fz��ؗ��:���j����T�a!�{=~�Xv���Q��Q�:�?�U�L9���l�t��5xl�lJ���ۭ�6�Vi��M�;�������]e�8�L0<��~\���6��Al㏤��t�,��9��_�u��`r�Sa�*���7r����G�[��5��i�\�����ɪN6���;Jcm�_����q=��۸�Y]��D��5J?�Wڅ��( �|�lhi��0޴	1�K�xL=���
���	�i,q�삦 mɇ�gPM�����C���FR�Ó���A� %�6���n6	LP���`h�h���)X�v>{1���3��Z���γK��3������q�#�D9��'�1��G���~���[0B�-d�׼�-_�3O`4�&�����0��0 ,�,�ґ��Z��cTG�)��,����~'Ns�x1��������ԗp�G|�H���5�|_����	��z�3�全���U�1jE��N�;[� ��'ܩh�!��N#�aa�7/ln��q]5��)����H�z2�KE���:��_%���bI�N$�4�((n��7�W�@�U'���Gl��1w��h+A������g7���pg�i�$�v�v�ߤ� �I��|t��)��	�=�&*�*��W���3��cL@�I�A�?jk��{8�L)E��K;Y���"N��@���1�d����� ��![�u}��&@jv���w�=[wY-����Iϱ(��#�1�L�O�Mw�0Q<����_�K-�I�)ki��>���"�\���߼P9"H0W+Ϛ�I`�4���i��)�� mp�bN��W1���y�cٯ�ϐgu"����M��~�˒<��_��`=!��H�2�=�s�.#3�f��E�QޯeaM�������d5��\�Ǿ������[Y�x�/��[� ������[���$�K[�،҆o�O�{vM�dZ�X/���5!"�2��	_� �a��YQЃ�=�]�4�l% ��A(��+ȿ�o',�\����M��� l-�p-Ξw�3�(#������-�99�.�9�h�z�)�Թc�5���'���L	W��r�u��ON�U�@	g��}�V*L{�m�^����_r�/9����f!$I��� 9+��M��L-�469�$����A��ڟlz��/V <NǍ�#x�� �x�7�ݼ����E��l:�:`)OQ~d	���׃~��}P;� �*m��~4E9�W� �T1G���f���l���#�7�w�Sir�+N�,X�	�]�=5ʄ/b^�ľg�J?U�{�v�ɕU��_s](Hz^��b�
��[R�F��2?�$I�[B@��Y�k\���,�� j?m��ې�M�;����י�zX�6�j���g���+�4x�G�?�6��j��J��T
��"�&ـ ��V��bI���:��ȷ����0<�\� �w:gG�	NM��=>I�kDt"��C���vv��}J^Er�����<�}9��i1�#BS�Ӂ~|U�9�+���yؐ>���)l��C4�Ѕ$<�J�j�z@x���M5�n.��z?��ͪg�#s%���il�E�?l02Q�K�i�ۻ��j��
�x�YC��J*ϧ��#���Q5���ٙ��O�g�x7~BRׄ�t� #��ݚ�Ų2͕Ѭgl�mn����]�k�^���
`�0�t3��Iv� �8o����z1/���cm^�8g ���Q�A�8����$x7��iO9��������-w �X��@܌]���G�gÒscبctXO~d�w�<�p8�	vj��\ݷ�6�
��Gr�<�0���Q��ϒ�0��K�_u�<�V����8W�q�C�0�����y�LihO;'����U8�i�CW	&z�ǈ�%��ʟ�L�E���{t�ټ;�k0��vP���R%��Y�y�\���bAj�i�_�;�RVFa���s�B�2g�[3�=�5$".�I;��a��s�� �c_��x	��1_1q���ݓ��M�b�ׄ���fv+�<`ڷ�8�|?�����������`��:?�Wĩ�P�׺���f�y���?>��,���z]��γ}��։����Bf����FO���9�� ������"@����������"
��5���h��L+d��Z���2U��i�!�0������&�2���������"3�8���W���5�S~�wa�X�V��U�*�j9u�sZ������Ƈ���B_��T�VM6D�ō�K�<a���']7��t�7/�;gm-"�㹚`����`w?W�3�O��I�|v����Q��510���A+ ��V�ن�ĵv�Hy��Pi6Et�Q'�@� �{,m04 ���*��Z�3�z�"P�|@C r˿��w�5�P>9� C�Y� LH`!���&t���NN-/�`�?Q��6���959��3	�s�<ˏ���e��(6�+��=�*w��N�[@z��z�m]6�7H_�.,� 
�*�7�t�����M�]f��$�F�3����$Q���o҂ߵl	՜�uj%?��%Ym�������a�x��q�T]�c_߱�"8WA�_��!e*况ʙ�cr���ܗ�s��z��~ٛ��ZGt��N��4�N��Ka@T��AL���$�� �>�0�L�8	8�|S��F�޻��FG��ޛ4p&�Pv~6�6[��s���[�҄p�2.a�AŪ�P	�����T�e���֜0x��~��[�tK��q��(,��x�f2VB��n����H�7��J��D�=�s5ǹ��\'���/o!�j���P-��²]�,�#���(�嚡{���u�͊�w��i��^um��'��}¯���`��+L,y��Fd쇖q ����xiT[*�����/�%Hp�Kvp��y��\�욆�����:�WgI�>vjl�b�\.ѡ�A=ʁ�I.��o�`�D�Ŝ}<LB߰� ��4-��QcuY����M��^o������T�SY�����i���#h��g1S�3��c�z��bU�'��F���$��Q+�F����͞���5��Uh�(�s�^cG�(�����>7;���%�+��N�Ԡ�8��&�H䣜��y��r$E �<L&��Ʋ��ٕ���j�W�$�x=�
�\E��A@"�`7��wIO.�q�
��
�y��t�v¼}�G�o��0[w&�^0P�j<���W�I���p�Q8�?ڴ�D�Oූ�?3���W�da�H�m�O�@���C3zL�nnA�wu�u%��[��;ܫC6xk��~�'/[����ނ�k$�U-������߱$,���b�J��	$������)����"�Y ��m{?��J�bN���MaD��S�K	NEF�����g��4�`xr�sBt~<�
7m>"i2���s���d�+�W�'-���$*0�Q54����Xٿ�wz�<��Lt�����K�:���nT����+���!�J�G{rғC:��v��':	VR��D�'���|��M)�zR�\�T��먞:�nV�(��8�͝	)8;��`����4c�2���K�w��rL��JGfO�^�^�\�,T��~�V|0��3;Y�|���]`�2YP-t�'��@@*���>75�_��OH�7�L�Fv���%���0��k�b�O�����b�HC���~7%G�}�c)����{rwк�s�u�����=^��d!x������ei�~ȧ����+���b�{�+b+�����ү�igL�_ܩ1R��^2�e���|F��h�.�`�
$�,N�#��R���n�;�;hq