XlxV64EB    8586    1820�~���)�k�<����'Aqk����7B&�j��TLx��2Zq&�;4�\�M�g
���.��*�A<n3#��\��e4��d�G�nΕ�ˌ��P�q�)��g��>+T�$����9ok�0���[8`?���er*!��:@��t�nj#�vͿ"1R�ٝ�����YZk��������euXy����*����O
Lo�ޯY���1{<t��ht�[��C��������{(�L[���t�:��[E6�M�b�� �]������c�,FD�/-n�<ܱ�ʋ����y�ҙ�
`)��nc��e'���{����<�@$�T�#�nA�d��l�}K��ȝF�J+�H0��@2b^YkHn�2�#[�;qBw;���B�O`��/�)弍����'�d����_軁I��J�{���f )�����l����cD�v�C���_�^>j�|=�ڊq
��8f-��ێܝqHdȘ�3@�eh��u�҅}�V&��#
�Li�e��(�.jnM��A�0Rc�w�o���>�;`r�`�Q��'��Q'ǻ�`����&5�-�Y��5*ۦ5dIǳ���I�D8���$p���Ɇ�O;;��0���3LL��N落��>J�>�nHv���1�5��x3y$����}�O���ς������k�+ub��*x�Ƚ޹2�ϸ]%��T���ן6g� ����z�s��v]g�Q)�bQ�
�1	���VW��K0��)�7M��(%��"�D^�U�Ux%��U�� U쁵�S��~�=�8̠���^ODd��Sz��QU�u��.o*�RO{�?Ô_�Ť��u�F��\�Ri���)�D�,�c6,����?�h��M�:0L݇�F�!���ʷ~ұ�U�jn��i�7�H;�uUc[�2�8�bj�K 3U�c�X|�0��ݶ���H)��m�O��`�:���R 1*K�n�PJ�=#��#<�IH���&b|�4@E���zgFԆ|�j�< ں�z+Cx�;A#ݰ�������FA\����
�cb�Ʌ�:U�����:l�J��{"���U�ԕ�Z�8I�cB&ncs�N��15*{�����f���ͅrZ���fU���C����0������i*��E��S�2���{��+�J���� �<o��.	f 7��/UvU�_;���=$�z0������g�et�}�6Q񅞟�5�;/z�ي���s���=�3D蠊��g�Hs��yh�V獓sg�[֘T���pL%�ӟ(���uc���X��C�ϳ��>� ��e��`���o�\L����}1D��*
�m�,�Z@lCZ�ö��.�ݵ�iݒ\ ANX�9�*m���܏��>�����:E�����JL'	�;�0R�þ�B�cuԩt��@����������۶��7���]l���R�`E&�\q����L�l���QD�u�!W��z�? 7`��	�ѧ+Ս�	.wBM�S�KtWc:�P}�D���<L�Up���uP㾥%��"�������v�#����BI���NQ��l!��}J�v^�_����e��4��o��C��^�l�\B�z�k�x�2w�\F�!�(5�G7��]��տ7�m[09'�3�4sSa�HXwF�=)WOʰ��4X^P�'�A��<�B}DZE-��N� jk�n�,�����z=1����q�2U�G� �Ir|4Q�+ZD�KC�if_�Z�����"#!O�wG$5.)0%���bG��q�6�{�W �Km�dG�{ȹNrE��Os�	��	���g��PL��G����e�\�Xh�g��x�U0h�_��B����d��[�lH�+�3%T鮛x�nec�eЛ�?B���]��ý��õ�8���I�����-�����,z6r��.��E_aٺY�/`+�:W�%�����
��'��*��l^t{���K��%'�(#�"���h���k��1���xv� ���
��'}&5�D���c~�EP8�����sn��|;l�xY�7Y�'�Q�M�R���*�E̫�s���{@�����b����Sv=�eT��VzE�}ʸ��Xkm�u�%��pzM�Ts�aw=N�4i��>DEH.�Ӯ���%Ǒ��˕�*}7)m7��'/S����@�O
:'	=z�3	�,>Fѻ��ɤm
�bt%�&1�9q��q���+�MϠNy96
�������<�hCV%��"�H�w
Sq��ef���Y�m*��'��?�]�8�)I�m��U�eH*#�5<}^�̼O�h�r�
��T���0��� ��T~����]����;��������5'�2���Ȧ�S���S']+@bo��ך���c�9C�a6�ƺ��y����/���Щ>�P��u����7�ց=��}ޟY��Ak��7�N��J�CtX���"	u~���n���c7��ܳ��WT�lA�)��m�����3�CǑ 3'��o���!�+�c �n����.�����A��U�&�M^F�b��T��:�Ȃ8vb���ytN�W,cVjr�v����̎X�Qꋻ�}��ҵ������7��@ǃkdμS��kdmsm���n�JW>�Ob��2'��|���H�V<?���՛.��-�+�zp�O���Å��G�Ō+.%�4p�-��C��U�����Y����.�b������Ұ��:�_�U���bQ%�Ɔ���|_*��W���镰���1Z��L��4�\瘐p ��_2��-L��eY$@ta�2i�5�^����Z٬`�
��,X)C�F+���+����X�~�����Ԑ&������U��/oz�㴼��F������+O���đ�:v�ׁZ�nm*_���a��PgUc�a,�����4p�!�ܓ��Q��/��AKrE�@��gz�����0�k��P�!a�.,�n��[���~�x�cU=�]�c&� ��̒F��4/K8�ó���t_��n� �]ꇃ�h��ƭ�	�(�J�/���l�uGpګ�r�Ͽ!����j�ҝX��wT^� {b�r�Q��������D�j[G=�-���ic�nҢ��%�i��TRF�c����@�i
���q��8$��&8�V�y��-�Dw�A���6 P\/@��܉!6j~��#J���:|85���<�c��	|	��S��f/��;`V�촻ҝL���S�| kVrs�Ci�*M����,�}?5���[�,��5�>��{��i�k�v�{#أ�W������{�&�4��ix�}x^�R��L����V-�<<��'�Q��h�c�_�BY>?�d��!$Q�H�|>�nכ�
����_�rP�[11:���)`��D�?���Xq��������w�X*π��i���	昆^����n�4�ϑ���o{��ґ#��>G�̗��Mހ7tJ2L�4�4F���p�����_Lr�3�1�f�GW�[׃H��_�-S�	�M8E�JM���}�Ǆ��JLY5�hiq��!Lg����H�/4=I¿��9��T�q8�O����T e9��L�"N�=jX��]N:�>G�@UE
?Yu3�;�m]���atim~������e}�CҔ��|��an������:�2�MKQ�6�����\btO�� ����E$��H2��'�ވ�9s�O�/ǳ�����u����%�u�Ɨ�+���U,�&V8.�
,�1�_#��ݣ'`DXs���sy@Ȑ��b��/���o���m_�}�&�& ��'�Y5�`ic����L��x4a*��&h��At#�"�}��z�X����TV�K�<nWփ��fq��w�1њ{G�{��I��ӣ��gȖ�7g�=(�`���L��-�1���󴬳6At�?U��E��r�!�t�V��_W���������3�Q]��+�:q������PPD��N��"7j�\	I��1KݺӁ�S��G��=Ɛ��2�(�y��؞���v�����N��]��*zY���ɇh\	X�~��	
6 *��Gײ�=4)�kU�"����z6���5���l-|���B�(B��/��O����j��Ʈ�%f�R�׻���R��t���N�C��!�$���r��`�Dc򷟤+V�4E��p�="q��Ԗ�Rߨ�\�T�����H���5�m_�V�u���F$,����ǔ�w�q���,��ٵjxMi�
�f
IK�R��3��zģ>i�U�9�g���u��{Ѣ|� �x�?5 ]�!�$	%�be��n�]�(h��` ��t�&e���ȳ�l�=7�^?��=��b��u�S��*2��"
D����������p��@�J�{���-sp���ir����}Q�֙�P"LP&�y���(mE䝮�.�^���d}��g��I��k0畴��j��-�(��0û ��y�o���\�*1A����@�`~0��z���s�DR����\�jf�g�^2�4���];|�D�|�����Y?܈~o��������V�VT��:��ŕ����ƓZWV��E��=^w�(ާ"5Xi��z]FA^�~�*]Y]��0�/��Ƞ;�y��Z|��J�L�Lq�vsq�ˡ��`�$����j�E�LYg;AN�i�w=y�t�����)� J��^ynI�=>�~C�� v�|���D\�߰�p7!�l��I�}��˿����ե�4=S�2N��j=&���3��xdCD��*�9y�H:�o��r��ܨ1PR�ܔU�����~#0��~�]��A����� ;iM�x�NI�!�R�d*q^g���}�d�
E��u��d_����Z�6�"�^�S򻗸�)W���EE�#����#M�F��`�QD�Ϭ6�Fvu�[z���XHzaՕ�u�3v��[�N*��x�N`�]�;�2b�Q�S�Dm[yU1֙�c�Z�jD��m��W���F�F��,�D3�w���WS�R�ikO6���Rf��xq�U��~E~�ǭ#����A#xY��N��]���3Ԓ��"-��\3�αJ��>
E�s�0ش�.,�-��[
�����o�wX�:���u�d�᥷Os�����n��5Ώ��&<�mq��͒�p���Ǿ}�4G;}VG&���#iy��k�bB�i�Π W�@��1(����	�5�������:�ffK�7MնC~0�T����x����#<�4�xݮ���0��k6g����=�yF�cه:$�y�Ri^�[kStgå��@�S�|w{�k�P��#�E������O��Au��]W��n�_`�:H�px�/]��S�D�N��ݿ���TǄ���h�BS�\9�4�k(������T]��:�:e�'d@�OQ�2D���z���T��G���]v��m��(9�=�ڑ�y&cl�+öu���p���f��ʟ�� Q}PXA��JX�!��ډ'�f��&B.�׸�����6.C�n�OG�3B�\6���Q�x�;]V�8o�53: =��pI�d���օE��}�3���i�����ƴ{�wS�;͋�/�۾ັ�-�C*�Γ�e�|QԮ6�W�&��x�a�xpo������3qeZ6';:���� _�ǭa�\Oe�<��xY�UP�ETJ��keN�`��Dm�l� �1�k���WFz�\�/�������2(����|��)�i�j|!}��%�g���|Mߜ����q6��¸΁�0�3hM:�O�4�s�&�lu!��{�)H�GDL�oQE�vm�t���y7I��#fP*��"Ϫ$q�y��r���L̐��د�(�X���/�ٸ�Ͳ ��H_�����ʙU*5�Z��Ǐ����r�\� ��|x-������:���#`��4:��H )�e'5�{������ͧǯ��QW0�q�������tq)�p�.F\x��� W�S�)!�#���	6�)�S�(8mZ)�tc8�5����������W�p�S���7�����c;i��)ژku�S�q��Ѫq�CL�h�A:uR�mc���;�=�@M���<��>�1��|�