XlxV64EB    2710     b70�.U)Qp�iD4pVCu����D��9�4���Sғ�{ �WGB=�rv�x��7g�l0��h�v
!Bd��O{s�Kj�����7ZO� Q�-�e�������v<��t��.�z<d�5���N�'��ϸ�_DB�7D
���y�ׇ�R��vr+���9�)� ���m�x"I,�M���&�aH,�f����N�m����J����1���ޅY��L���y$&Q�U:�|���u��k�X_���Z�+m���uJΟ��Q��~c��q#�s�0P������8v+��*�<.��d��S����/�N��3�[���|�x�S�)7�g#��JH>��͒`�*n])b�:�e������#`��h�.!bHAe�h�,F1����=;&,��iV㭥���7	+�Ňθ�EE�Ԡp��	wַbxp���u���QE'1��6ϑ�B�1��Q�o\�|'���3<���O�^T�QҔ�R-mC�l��z��OH�D�E
g�X����}��y>� 2�AM~W���m&��k���c^�`��3��9�!,Y�)��@Dl�^`4�d�u���w�6)l�����=������,Z=r��
	H)]4,��
�@�Z߆ő{���2���`B���d���K����F�)[���G?��R����0֙w�\=����q�
08Gc^����J�T��)�=�L�}����:�B�u6�&c9����.���o
4'==�����H��jD܎�A�H���%���:��ؔϏ��0��Z������IC�>���~.;�6:p���4_䷝�X*�R�2���u ����Ⱦg�&�,�f<h�����.k�T��w9v�NRÔ�"��	�����4=�g	�M0��%�C�į.oB����t�Ma�N��_��O
G�9�a��.��U糿Ԍ<�NHRٴq�����tb�/9A�����¦G��C-��;���p�F�;@��~<wR-�S��o.�+<��t,�s	q��b�cY*��3~Q�z� ����r��kQ�K@��v������آ6�a�$:��M�2�+]5N @I;!7KmR)�d'���5 b����-m�֜�����P�H����/��6���@�X��!���0�Zv�0�Y,��F�1Ml��1Z_����FW�'��1HM=�p_�AV1m�8�݆yĚ�cL��Y	�|��n�e�[�X�ʼC]<̧��IXJBwp��
�ѭ)���Z�XM���R��R~��Xn��(�3���"A,u��Ɉ3/3G.�ŜZ~�}h�g��$�_R��ގI@n1y�n�Lg�,&9o�@�5��/�[Rي�\�oծX���?���Ӌ��C.�m�:�TR�8<v�PbS�22)��� ]zn���U�����~:�f%�Qz���&�&O�:��W�lS�ވ;����
<�W���$�FnM��L��8�H������9��+����ڣ��K�-�62}����t��Jpǩ������uR�h[c�#i`ۺ�jqx�fM���O�'9N�"�`��_fcN!B�
�ډ����h7�l}La��{ r������@Z� �5�i�\NA�h
3�*�0p�[x�-��8�Q�R>��/}	�฼�i����پX����� K�qW�l6��m(\�n����U�Z�ۏ��̳$Y��m_X&"a@7֖=aH:��+�Y�V#��Q���-KQ�@���1�=�i??"z/� cL�m��.�}��}����֜`���բcK��bUKPR�f�a�c>�#�Z���f�h��Rkܣ$@l�!�۹�%=��t3=܊	��S�pi�iӦ͚�]K���r��䎠�l�o}M/�3��.����>pc�n`7�=H�k+��r'h��y?�V߯��@BЧH�Lm!��:��\$^W��f�LOi����a��]i�3`�3g��צ{$�A�	���	�rZ��kn:P{�	� �;$��uS�L���;֊"��5V���@��K����)s�0��%��򢅄�mxv"v�(u�uᆐ��َ,x�(ݗ�Q��T�Ԇg��O~p�V���µa�%kf%��:�d롴�ἲ�!�1�%��B{N�"ϵ����g �������݊?���{ֳ됺�kY�E �6)n�,��0���`T=nE��e�0��������l��9y�x ���v�]�?�f/�[��S��g6v���)'Q�v�����ySQB�#�s@Dr=��~�	�y��r�����;�Zԋw���F��$v�F�ˑV��Btg�}C�j�`�4�DT�z�JLr�0C�J뽒`b�-�K������o:����Z:���'����F��'�q���u��E?s��3"��]��V]� �Pt���$ܩt��|S;���q�b<Št�����Ӿѡ��cadszX�	/���z���C PAn��y/��@K����Z��	Es���L徏���/1*K���c��;�G=��i�l�lM�l1�:*��mթ(�-L��k�o��4���|8c���@m�~�D�s�ϴK�&֊���h��ͭ�{��mC�{�K��m��&����c@2�|�,�x�Ep#����F'�+K�����N R
ȓ 9�g
{���8�Ts�~�:�;��f��i����&i���aJ\./�X���ȕK�[q���M�%1����5�Ɏ'8����hWTo�)����#�����fO^�M����X�o�?���V���x�Cu逰D����_��+q�����>��.�_�[�Yec�D���M�%Y�T��y�b�A̪cI�W7�ǥ"	�j����	�U���<ޗe֥�gA�[��i���1�� d�"