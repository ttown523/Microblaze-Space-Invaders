XlxV64EB    159f     840"b��ҁXc�D�x�۽A$l�e}I��Y���E��_(����N��H�9�7l���+�J9���-:|ǙJTݭR��bP�/9sS�$���^A�v �Y���+�b�v	{�Vt�R�������Wc�N;�*G�`����@�s`�^P������� �]/�I���$��%2�t5�g#�*A�-�͇�^��HK_d���'C�gn������T�5���W���?g;,�s\�2���tm���v����֔��ԩ}�f�Θq��s0F_�t���>���˕h�L,
WJs�kf�mf�aǰ}��<���� _ȟ��1⺸�Xo�-�D�Œ�r�@]�#n4�޲���yJ]�='�!�?v�c�~^�Ft��ٖ�|���'�Y��av^�(	�%8z�Z���8�k~4��p���c����Ώ�w��X�����`,
R�������$M$�Ezu;�퐒3drN�,���Yѻ�G�^*b�%'��%�l�;�]+߆)@��s`��8N�U�Jv���&���
�✥�_�"�vXa����ñV���3�⒲�g�Q�q{uԫ:��3� �x�M�9�WD�C8�<U� � �vS����m��G�*�V��#����wۖ�����<n���-$F"	W�FJ-��}z��D_������8�o��f��ږ��nwO'0�˭��$���`�L����<1l�ѳ�0sH�CQ��S�\l5sC�])=�)���ɰ2�?Z��=0/'#�#!���jl�6q処vq]��ڭG<T75��U�d���	,SƵ��:LXL�d�fa0}�.`�7G���zR��X#w!
��GMȘ�A1̿�J��Ws��T/��z2[�_���h�]���.�%�x\����zz����V������D�?U�d�藿�4�����d��g;��Y�i�WM<��@]O��3/γ�9��_pu�d�BM�r�2��a|Ѵ6�l�1J�}z����!����j�fm$#3k{8�s{��D�y.:�C��� 1fD�^��������ŝ���
�>.q=��)\-��d����#-��q#z֔�?�:�u�q�	�������
��d<fP4%N	�������Z�u/#�3��[�����暶�lml)�]-�B���y�W�����E���BJ㥏x5�EG�������u>F�~v�34�2��["A��@�)���LW��i^�AB��x���l����ϒ��G�;G��ſ"9$Fr;���Ī7'�i�s���Ŧ;�Ac���8t���a���՞M���#�s��3�!�Ȼ�9�^|X�d�B�>��r�_.X�U�m+@鸕*��P!{@%X#R��G<N�R'k����a*�ZdZ�/2<���.��'�4�W�6���Qj��vA�.Jh.�㛂zN��U�c) �����xJ9���}��Ԡ�a�L�qM�F�8z !ϓ���*~�}jr�z�r��r�Jڜ��d/���a�������4��Yl\?�;����Tۤ�]t�a���_�L~ 9?M|\�ёF]�i��zv��brZ%Z�{�@���P������f��=�x����@��qj�K���HG\ģ��O��ȁ#���|7ҺPA��[���
�����HEs�M�h$��$��7�1#��N�`[:)z]El+� �d�@s��� q3�J�R�0&�wr5G}�g���+R!��L�1�8>CL��7G2�fL��Š{�Ž�"Phw���+�M��<�_[T�K�
m봞t���7b	0)O'9��2}��W���Me�Xo�i-���gz��id*�r�Qɔ�Q��̪M�x��?
:ƽ�o�d�!�ץn����p���H;���_��8e��k�Gz�4JA����ʡS5���(X�]�!�I�N��K�y����p�Q�>{S<AЁ��"�]<��o�R;ASS��w�B��Tn�g�w���V,-ʕ�	a�iH����
��q[P��V�[|��d�F=U,�ُ~#��2�9��qfBK*�q���1��iF��x��q![���Qh;��n���4V M=��|� '!��]"-�m