XlxV64EB    20e1     b40k�s��̸I6��M|�����p�*P�\�~�$�+;�_^רL��,����$������}�C+}=�Q0_M�'VQX���4M��E��Á�-���2��~ӂ
r[�b��q��:j�vp�w��@|��E(l8����r�w�B��A�6q�[+����/v�n�~e�w=�8������R��1��\�,���!Ԝ`���-��Y~�t�K"��]u@ȹ,K��������5U���SN��o�o�He�'�q��f�?�6�)�.����?����3N�ZlҬC��7M�6�=���θ�"��ծ��y�Ǳ���R7h�� @L������ٮ��&і���]��A}�6Y�%I�0"-����O����� �[g������ ?��|szu��w��N��+� �R���[J����M�����I�+ӞyհYA:�f{+��bb�m�KV��N���U"T#m_�($�rT9ʰT�3���4�ÿ��N����	�a4��15z�+o�X����` ^j�5���� x�_K��G�&�`ř��Yk��:��f^�֐��)-�~��@հ.m��`��?�m�%ķY�'��/���M�rI��9�]1��W�O:k�"�I
��n.9�b�X�@��?���R�2ՁL+ȧ��V�-����D	�))1�¯�"m�W_���� �5�{�$G�NQ`���玙`Trq�y�9���K'L�N�<�[�u���d4� i��"JKH	���'�Jm�8��9�O�Bg6����	 v-���h8����쮏������2�716��g=l�Bb�徭G,��k�N�����eD3�F��ka��6�3���e°&w[k�Iy�5��P$�Ahy�!���
&+F
��J#a���E�Tq��
�ZN)�
�O�%}c>S0"Z�w?�Ђ%n~
UB
C1�W�}�.�*�JĲ��5�ۛ�V�.}�ddM��K�:��J����D�iA�5M{��ȅ���
�
T�3�+fYT���Zs�:�#��J�/O�h��b��[��v��vg�r������n�/�9�^e]���A�;=��p̧s�sw]���m!O�S�O�\��2����3����\-�Q�E-&N3Vz����y����M*ͭ"8$���h�>���!�h�v�:�%�j��c�U��eb���
�0^��p���Z1��҇���9<�(��5��Ptgz�k�~>r�_��"�����>�m��@�t	ܳ�w=z�� }!������3�"��Q2 OU�+5�c����^���[�/.� ���Qq���K��<�J%�liۧc�š�Ey�fh��bĕ؁��AWqj7������c�Z�#3*���Ӯ�B�ېG`!@�{	�2?5]�|lQ� ���p_>�%~r�o�I�G�}!Ia!۔�F�����;9�����kJ� D&{�L�����d�B�5�JM��s#D9=o��߂��lw�i2��$߼eϞ_U��NxK�{�jKv���@�?P�YU�Mb՜���W���ڌ ��>d�J'�a�_��(��ZN#��$�z?d��3��r>���۽
L0/�+&���rR��K�	��h�=隱�z=5�{O�y?��������"�+B��o���u7u�`�����4J��3{��Q:�>��c}��vkv �t�0Ug������d��t����JzW{Q��c�& ������#P��K�s���k�[��څ�c��_aؾ�V�a�k�wj���X70��nbY�`}E�NƝ����5����in��V�>R��������\��A���u���Q�U��x��v��V���H����. x���+WM��ӿ����1 Sw$�T63��w���o���v�8ET��qu~U;P��h&Uc!g�@�z�*0!��Ӗ:������s��
�Rx	���*��v��n4e=�(��<Hӊ�m��(���%��E�{�f��l��	�h=��G=�;��e�9���4sp1�WȯNM��z(`0ݹ�4�ט"�-r����3�����N��7,�J�����}��|�Dw���MKݳ��s>�F�~}Χi��/����}b��-�3[���G��� ��#ƙ���P��	X�v ����B$(���ñ��n�n�Bv�g�����R4�>e[�{3M���U}s��5��;�&ơ�6,\K�2�4|V	z�p�z�N�k��&mJ�WO��9Š���}�9fX&�t208��~f�?޺EK�ip�_��}W���;K*�<~{�Z\�.�:�V9?��ysA�x���9I�k�ʠ]�1���;�]'L�J��$2X4����kckh�F�Nq2u�u��� rOAM���r�g� �rGE5��K h�Y�&��u�K�In�_ 1$G����|��ъ��z=��&qe�.�/�r��������@���=>fZdجl
��\1N������m���|"���5(���oG�p^~��8���É�k��۳��׻�q�.L�ú�$hLy�!Ni����������Q���W�H&*0�B�?oE;�oy��-��ͅ�#�C��u���E��B(Έ(u�H}�,N:�aEU=iK�R�5�\�L(_�ggn�Ris_ո^#�������鱎BPy�,*�������
 �|B�k{V�@�}�^��~����SN_U� ��ڊ[zA�lR�\C���U>����{c\ey~2�Aqp0VnF�v�2��${�,��FZ�ȏh_��0k����d���B	z���i�]������� ��}9�����^7�