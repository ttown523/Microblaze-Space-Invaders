XlxV64EB    2aec     d10���4�A�� � �_�����b"�k������eV��ғER�{�:*KM>���4����<�ׂЮ�'�B�mXCл�57�ad�	XJL���0m������,��-�>�(���,���U4B�Q�9m%�������'�78s�ؒA���[+^J�cƁi|a�!��Ğ�nܩŒ2�F��%���$����8�0C�L�>�U�׋)�s2���	U}"t/e��l��^�d�J�����*!�y�F��jW8�=�X��I����}�#���WQ��2��m,'o�TZ����]�*W^1�'��ĔX_���(n��P�Q�����)��2`U��a���I�ׅ`5X���S��F��ļU2�+n�Z_�f����x%\R Flw��4\�m��`t���h�H\6:��Q�`��q�ppȘT�o۾'b%#\jD�dT9�
$x�q�ǅz������f#��kʦ�I��N�&~6.�^:'w���S��*�ꏎ����c�����ӿQp8w��9V�6lM���ø�����VI�n��D�� ��8XӵƱ8<&�f>B1�{{1�G�������pA�֎{�{�0���&�/�	q6���>����{k?�mPQ��L������R�:<ğ�;c�2y��
�L�|T`lH&:���c1J�W\���&�qu�BN�C��f�u��3_$���?y~]������
l,Z�)�C�������v�iIx�x�M"��}4�b0��;�j�9���m��!�o �
��{u8b$���J�^�'�c�/@��6M��4��gٹ����7�ߎ�i�_<��TAk��M����S�^�d#Hͭ�r�������Bq3�=�� ��mS�*�t�]���Hc�Ȫ.\)v�1X;�g��qd��(ƻ!�����;�$ ��5��TI,+]b+��*�Ya��w��i���*�<�x�H�M�W�-��]�$��WǸ�E����w1I#i��[��s�ʔ����MK�*�BVcN��/�e�c��`� !��Z��o���)�zϖ���.T��Mv�,q�t����4�&�$���['D(X�G)���p3�uv��h[���t���7zZ�(�h���z��O�`�n���+:l���Q�Ք��_�ev�������J1a���D�?���1����L�y(,
̗���W�K(�<Up�+�ygyu�=<�j<��+�)Q(�*�P-�8'�X��<\��|E�܇�6������Ǖ?���`���Ԓ�cБsW�\x�Gr�x;P뾳���W7ΏE��<�q����s�u��'�R�2�7�/�����p��;�BU"�x��T�|ssm0�n��%/dڥ5�	����"y^�I��ڱa\��HB�	��zD�b�:�U�� +����3�Fσ.��q�۰�I	�e|�K�6<�i׏�=��w�UsC�0������YRo��q���Ơ+��a��M7��0�4�Dt��"��A[�3���o'q�a%(+��X��O��l5k|���#�n�J�ڈk�T��WM�D�L$Bm�f\�I�b�����T6��觹�I��b��s�8���#��Lɹ�l�ޱQ,5�OwM"03b�3��؇}�^���>��C-<K��&�u�8h���*]�R�(�_���Kxe8�ucf�E<����l���\������nåW&-�z�)q�cR�5P��n&|��ʣ,�&�몣1Kʩ�]�v\3��\��.��\��f!��P6��e����>8���oϗ�L�⫡�MKY8�K������s0�����fv� ��5䱁�JB�j +h^�ʎ�K��.�},}���q3��2A �����n\�CO��ժ#�x��ՙ`�[�w��]/&���LC%�i�b���G=+
��it�?�n�T֫����G�]��d�ξ����'@�������a2�Y�/4�B3��]hIq��awb�P�߰�T��"b���}�W��A>�g�~\����*�c�[�>��\�#k��6�*�HA,��M��óE�M?���^���j}�z5I���������������k��6�EDs��4��`�R�a���YQ��e�t�\�I��`��Ԝ�"���I���.%��,j���̍��!��:�5SZ�=�.Y_IQ�=�C�{Ə�p(���'X�t?j��'3��R�p���me���@�%� ����C�@CEBh�7��kʴ��bK���Q��	������b,��@"��

Bv��Sԁ���0 ��Z�%����E�������Eݬ.o�D��	�+q>�!P̵���*�x|�i�~'!��?�DI~�ٺ���.��wk��WNi���.������q�/M�<!_�)�c��N�?�S~be�[�G�<j���f�o}�d��+�r�깞����S��3G����A<9������4��F�v��dj#�G�h�m[�,�d5F��)w�a<|�T�O�*�
ߥ�v�y2U)~��Pb���|�aM�&a��wZsD�������{���{����''�J�%�K�~)r��e�) �������|v�0�+�vzt�/�M�(e�B�ۈ#��R��=\H'��z�������)d����u|S�&_z����g�X��D��,��?o��J���,_�
h��vZض�;;�����-��>���dř��<0vN�#10t�"�VK�Ƃ[�)�V QQ��7��BXS0be�!a.����p��==D��4un�����u���?S�cm��{;�@�Nt�y#�/g,��$�����_[�ګ��\Lʤ�d*y��q�r"n�㸼���wYO���|�+	��%���g��Y,[FU&&�<��;8�K�7N����T�r�q�� �0�=d ��T�8񚌋M5�'���g�����"�4�X͐7�ǚu�i�cm���>�J�%G3�ʈh����̚M�Q��1���1fa�ϣ��쳢c�i�����7����z��A��g��<��K�񆸺/���,#q�+b��2͆iѫ
���U}����=�h/\ ��Z3��^��_����x��,�AQ���y8Nj��@=���y�Dy�y���7�V�a�x�iC:�Uf�W�>�7���}�F��\� ?@���:�> �k��|�||��@�8;��C�R��%�� 3�P����(��z�(���������E���<l�$<��uoQl'��rX�l��(�,�I��(:@����y<�x+'����&SR>�15�kVV��jO@�.