XlxV64EB    54cc    1000[�
����
�0���8�Z�=y�\���G<w���SC�=71(�6�@����Z�b�g����`�fc�>ȣ��z8���?9� �~F�P�������<�Q�fra��ف9��&�e����p������Xt�y�f�pZ�v�RI�|1?jvi��GF��?�����X��Zs�~!�?�}�(�����ޠ\\ʨ�n��f�h~ߋ?�|�g.o��� ��r�t��v43ʭ03�u��.�f�J �d�ÐC�(M���fv;���f�#,-x�����ˢ.^;kJ�.K��E�����M�R�D���П�&��Ɖ<&I��_Y<ָ�UK�2KT��`Ȋ��ra-X�G�>�C0`�iW�2�|�Y�؁0���G���.��z;�I̴G@r1$+ƈ{Q��m�o����<�rMCݖ��Z� ���q�פ�4ܭ�;�(^�ĐF�miBg�I��	z.�-���VDYe��b���
d{�oՖ�柗�Ӗ��Ở�]>u�2`a�cv@�SG���Bf�f�k
���O�Zӎr�Ox����$�v�]|H�\	��k�bb��K%yId��^�"���LY��8�O���GJ��2�0�T'�q<�.ܛ�:�a�&(� ��ֳ0)-m�;Q�>43�x�*�yP;�A�Ҕ`!cێ����D�|�Q���~�m��-�M&�.�Y³Kz��e�'��� �+,�x8������l8i��<�b]�+0b��Q����^
��.E�`?W�y"��՚�5�	PXq�M(��i�"�G7~�S�t@%uC.XD�bH\�V�u7tN^�]LÙ��y����Y<��6s,����uة�3�&6��J���\��s6_4��V�@�gKVP����<S+�|�L��3���ٻĽ7b�y��9 �KYf�m�C�N1��ZF��R3���KY��Nc�c�Jh��a�D>kn�%[��*�� �1�K�/[��3܌���)t��ѣv�2�C�q��n��X�ԭB=�R�io�(�GV(d�_M�zX��+���l�.d?�|ƽ��p�O6v�6jh5�T{�s;���>�@�s�.��z��z���r�y�h���'��n����17����;�z�?�Ma�L�I���J�L���nd;8�8�j�ɏS��(�֭��?7�����,�z�,|���Fc�a���e�2����@7�~C��<� `N����&Q��	 hH�m�lSTd\N.�3<o4��7w-J
M	)U\�D��'��D�%	��	�q��O���0��m���H��xD�ݮȀ(ON	�>�X��x?SmN��o���@��h�,n�����iS�˗�̀^�	q9[�x����G�b3�8�-�r`Th��O�ۥ�׫J(�b�;AG��Q����|j/!���P��Nu��J
"��n��`��3�dS�L�6��H���MQ>�`�/TҾ$�G��?���Ň�.��g6����Țq!�F�:(A?Z�X�z�h?rF��oC7bo0v�B�����h�OD���7�h���MRZ-V�:��5ף�q�'�a���4�r-�LA}w��i���Cx$��/��*���x�Yv�'+'L�x�h1{�56ƠD�T��ܫ���q/�&�][�n��T��vpW&���-zѦ�qc]Ɯ�G��X�(v��~\M�N;�����j��O.r��/h�6:N;czqM����ڏ/�ؙ���^�ʟ)�J�7����f��z�f;	��=��t#�e�T�M��Xq��g�?g'���m�Jq����l�����Y,%�p �~�da��U���i��(���c��vb��ת8��zz�Ylք��;�H�$(������Jc�~�B"��z��I��K=�����s8�Z�8G�	1K޿�	6j�2}�S�@�7/��E�B�&
�J��&����"�ū���j����kE~)��}�!@�{|�y+�z+o?�Q�Y]8^e��B1��b d8�,��D9䩾:n��P�����]=c4͡dt��kO)6�޲z�gz4�&�TsnI���'O�n��i���Ѷ��� �+��l�[-��If���XI\	8'h�h0i�ֻ|ʺp�|�8EY{.r���(�b5���ܭ^C-E n��!Q�R'��s���I�<���g�l�&�T�wsq~��2'|e]Ac!"`[1�I����d��9����S�.*ِ�о���xj
3�4.	�Y���v�tkl�M��m���%�F�_�խL���]��������;�.Y��7�ͪ8��j�_,U&� rd��?l����:�5�6mDa������L+xӖb�P���)���.�9���F�>.tHj��u�¨�y���P�w�q��_�.٪��|3=���\�CU-_^��#Ku�9�`W~,o�<'}���v�B���}�6�+N�5������Y��،'K�7���I���T=��p+<��&����U�`�������ޢc��0���U�vuye;O�yy��9g�1�X���%��Ty����T��;}���N�[�/��YF^��l��S$3��摕b���ܢ�;>�P �j	�9��Wբ�U��=�t�C;y�Jm,ʢn>��5��}�`���_�@���^�x���U��� �����ZP?��9^� �ex;]�ш6�s��b:�D�	G$(s�%8��:CÞ����&���*�R#��r�"���	��u��yi�6�}�b~bBz�;�j���m�|\]'B��4���n�*��3�K����Xq���W&0�{KA*��9�V#��������çX��3xIp\�H�Ю�a"�\���@M�"e�5�?��6��
^�X�� +��q/����\ٽ�o���h��Tl�o�)!��ɻ��?ɶ&a��=�;���ɬJ�`��]4��i���-Mw/B+��m/J����Zg-�w��}��DD�ǋ76�͒E~�D��؂����f�?0s�� /�6$/j#����.�����!y�;v��6z(E�rL�li8w�Zڹ�7��'*�h9�HbMk�l����/('��܊�N/Vf�û�}�f:7��$2Ԯ�4��Y�{e���I�r�$�]�K��Dܮ9:hE�x+PQ@-BT]}�W�r�E7�v�߫�4��ٿU�S9��{��)c���M�}"���Z02�2/n��O�]�mU�peK[���y�=��"�@�Kv��P��M�`a�R����j	Ƀ�9�\FV�I�,P�S��ï��7J84��<&�y�����:'�)C��G�4K]S���j�o�����uT��VI��S��H���#�]F��)M���Lt��2(��p6�M�~��Ssb�faLC �����#��#9�.��>�3�;��IQ硺E�0z��-�C��G��A��Dd۫�,Ǩ��|F0����Fl	�4�)��Qu�³�G`����Q3kW%��P�m�%0�1,@��T���t�B�/%�(��2¶�4:��T��D����.��H]s;b-边�!��*)A� )�-Jk}����h4\h�B<���s����K�I+�N},�)�a���I�z���'>d�^�h��m��Q8+�f�Z~�F�Y�MU/����\�)��0d��*����ۤ��Q���k\ GY
�Ѡ�ah���b[��������'���E$���VE��<Pۥ]��$JݗmP���J�==��"»|��&@��q��e��s���B�����_{��k�:?�ӱ�)�m�co&�E	�svG�z����R(���c`뚋Wr�����s�Tt�l��1��)0���"�XΧ����[����BE��z�u�B��3R���`,���[��he-�����D��չr�(�L>�^��h̥�X��p��G��M
+�.�'h���+����ӥz oD�E�O�銪���R�-a�P�G�u�ł ��!�KVv�-)�ro%=�Il6� 4��q.#�˂9����m�b��2��78���5d��؍sŧ{��4