XlxV64EB    17fc     9b0��b�O�� ��z���;#_1DC�B�����hN��W��R��\o�C�0%���C�E�2��_1d=�y�����RD�GKB��ż$I�J�R�^Fyp���x���R�2�;!�?��� �
�|�(���H2èW��ONm)�k�N���!�� I��u�e"�'�]A�TH���_|�E��7&�������0�����y����c�k"����eJ_��ኙ�^-"F"���jF����k呄�]2mq�,8ӝ��V�7;�2�Z��Y�a�uZ,r�L���ծ�+�6*=H�TB�{�|m�Ý�L@�����6;��_`W$;��Y��?Xv�/_xr���L�V�b�]�6��g��(}�,Vg�&݆���mE���s���Y����yh���_
�C �*�4�$��%����� �1ݚ!�����A^4A�K��rP��K�H ��=�B��$~��@�o0)�@؛~�zQA9HRؙ����Y��x�,�:}�"���I5�9;�Y�@H���^l��o~�]{1|ܫ4p��?0��]��?�e>1I�P7��t��d)��]�O���	�C�z;f}�ɖ��U�WV��MNk����O]���Ѫe"#AJ-�y��OT�u�CS��� ��,�f^�fJ1Xf-�*Sl��F/~j�f�I6J_��4w#�]��Y+=�KP��`N�V���/�d�x�D����Z�*	�|����.����^+�4^&ؚ�+&�nga㸘����N����*�L��#5~���_k8�̥D�/Y�h#�уW�3I$c���Ac���o�`�e�](8Й����(%i�ս���x��?̜M�+�xd@�/U���<�B,��Y��}�`�� @��{����Jՠ�xe�P�ύu���v4p_���!p��bǒ;�VA�/��.$.y'�Q��6`�PAɑ��~�o5p��mRǒ<�8	�Qj���JC�WL�ܣ\�3�]/-`��K���^��2����Í�"_w�0א��(6�� ��!�s��r��"�K���c%�, 	�Ԋ��K���_j!�1���*>��q|sh�50NSx��G�=�@8|�5��ċq&��{�Z�y��V�eD����9+Q=�,�����B`�-�򺸣3>
��������>?�镜������6,�k1�%
)�p��ȷ8%���5\��(F���Nhu��A�q������l�q�b��{�2�~=bnG �VlxS$ԏSo�L�/lL����_����s���-�zi�Ql,�r���É�5Fo�!��Ѩ82�'�K3�:1�0|�M�&�mhL��^]�g��J}�<a-V1���䤏�9%�ˆ��k
#�7;����B
es*�q����UI��O�h���*:�[Y�~�H�7F$&|���q�DI�ER�tg���zb����V�W��l]W�(�J��t��yV<��Y$���� psv;0�"q��������`V��͟���Y������N�<ֳs�9g<���:Hdd�޼��D}eSZ�����%
�"aY�N��a�_`��Z�$lQ�Ҹ�UR��c�i��uC��uW�'HD�5j-MyR��@��,�����A�Z
]
O�4'}�hg���|̏DY}�mv�L��24q��E�:b؁����3t�*��ׂQ�~j���:��5���c�f��:����}�CG�i�:<��e�N#&a�h����~���dd!U����Qn�Q�1j͗�Vd�9@f3���f����Љt7���{d7M�}�']P���"yN�#d�$����(4Sg|�B��	��ϓ xrΘ��@���@��vc��,q��ˏ?T#�au�D�^��=�π�)(�-ڱ��2��pM^�f�A�w@���pg�ؕA�`U�Lbt+�$POk��p�I=�UaD�8C�2��
iہ_���b�=mr��#}a�Y�+�!��ﻜ�,[����^B��z@W���|�p��cB�h�o�&���O��N�
hU�_����]e/�sb~��?�)-q�?��
�����2��g0Il@��~��~�WIӰ$9��lI�I��22B��+�$�[rǃ�kG��y�V�NM�T�g��X_�{L>	?�jF��A}�?�U�tHL��ɘ�k���m�2)�*q�x<�N�0u�#O�� ��anbJ�"J�j�_�fL�����Y�)��o����e�N�X�.�󾳚��HFq���������ct��MV�a��0#�+��מ�2���>�b��⼓\8+eJ��	2:7K|�ʼh{�CI q�._�A�Ғh6TP��"G�@���M0΁}���C�DX�8�--�=���C1����[�Z�z=�g���l=�L���ѩ����������m�w���������!�ȡ[j���*\R�_Gz ����-H�I��"�^Hk