XlxV64EB    4734    1240���P��բa�
��
��l���f�F��U$��e��21���?�OH�L'��6�r�|;Nt�ߺ�fו�NJdW�f����1�c���t�>�8���s�f!��1�%��*����:����q�ܘj"����5	�G���f�7n垄(JQg����p������M[@y#�h]Y�V����8�$�f��@�u嶇��d��4���m1��K��jjC�j�x[!<4�����J������� 9��lO
Ȼm2���$@D�#�H,_sG����}\��]\-�\}��X��˩�JΙ�t�Ʌ,���U��)�p�ځ������s�! n���U^� �=T�K8qYh��҄��ءOV�c�K],R� �Kܔ 6:����-x�O�����u�����e�A;�#�-�m<a<�W`���$���m��8D�R��T����#%TZ4���Kx.�s1�iOqo�����,a0������؜���"�W��f)/��z�ƅ�?���&/��+V���%O�y�\
�"�~���[��<��0w N*S�]�;d�� n�`=,o��n�"��GӞWp�o 
qO��ܴ'w4��ۅ��fW��+�	�fb	ŜM�b
��9'm������p+���I��-l=¨��]����ŉ��BF䤐�YQą�(D�\��)?�>y�Bj�+u4�c�$��:����L�C�Ե.�p�o�&����v�j���	fN�R�6-�d�(f�i�`�O����r�&,.�qr��������K,�(�V���~(�rä��|����)E0�ʪ���b��b��XQO��������%�*�0)O\+mQ�<ߩwM���l�NsŇ:� <�{e%5�huL8�ҵ��cZGz������R���bd�<h�z��'I���̒�c� "����/n��^ȳ�JMM_��]�{�3���1P��qg���j���C3���w�X9��ȳD���M:�_$X��U耻�Y�z�	��L�I�M��$��آDp�)��]A��muh)��t�@왞)+'&�n8n��=/�Љ8��-�m:��M��H�}AA�>w�B�C�'3]�0uĻ�j�l�霖Q�y�����=xo��<�Y�ߓ�C��e�b.?�IL:� 9.4q��=�[��]-�*���K�qf�3ȭ&�����:W��Z?��/�������S3u�J���B-�,;���GX���Z���d�.nO�#���Oc�r69o�(;L� v��vM����F���dP w�V��:�:���.�<Cl��ʨ���<z�90�p�Q50��	>�:~��*tڔS�p`��V�X��$��hE�"z(e�o((�y�<U� ��ьS��U�:�n�RK�4��	��	)m�
�G��D��H
$(��P����C����ތ�j)I������3D�K}Y�����[ �F{����鲏\��^=��-?c��X��u��,�oڭ���	]@�o5;F�5n��)�S���@4S�=�ߑW�wΗ4�S��}9�����iX���&���|����o���xR�C�\u<�T���c�C}�+��I�������R:|]��@��j�aB�w�M��y	"ȭy��^�}DiT4�mE(��5�L��[OV\1dЛCB���O���b;������3�r@7,ȴJj�\����5D�7�Z��{�v5^	ˋg�4� �����$>��ag4Ks	�AdǦ^��d�?/J2j��K������ (޵I�0��z Xl���@*ti��c�0�ɳS��hY����K�+�MZ6;�WJ�e�����?h����ӊ��?����t��Y>Vy��m��N ��MҀ���bT�%G�Oh�J�������.�XI6n�z��{:���fFެv$�G�Nf���8�'��Q��ѓQ4��n4���/��-���"�q-������h`����fG���&(�����\Ǻ�����I�(��vq/)U�US��p��C��,���v��Z�$��вe�����P�Z�|�1"����L�|t���p)~6j��Z��~��-i�'N�<��څY�CD��M��l��,�.���\�K7쿔x���R2�1d�v:֤���S�zЋ�!�� ܴ|g�pt����wϮ�/A�A�r�8Q��dxu鄛��e����e��B��A)�X7���-�a.�Ɂ|>�_p�%���9�!x{�,��#S.�.��f�$l�~�48שOw�j0x�ז��Whz����c.�\	�E�)�K�Y��������O#_��?��E;�k��^��G		������茡���-�������SY����|,~DSg^����V#��ʅ
��i��?���l�N�z,��<��F%"NÜ{�e�il����5Q>t�I�1�G�9��히�R�����!�s����1a>�P�>��Ӫ��r��nkq���_����W��B3q��a�Y LM�; E�{=n��$a�''�,��8x,���w��]���e<�^!�m)��~ql��ֽ�Թ��
�������v�����P3p\����|ͥ��e�M*0�Mt���)vK�� ����V�r���Z��}L�EJm�Q�b���: F���o���H�o_���u{F(��6��e���6 ,�g�͐�׶�|/�-d��������eH��'����>mB^��e�Y7L~���{sJ�/�\��c��1���Mp^
M5l;!p��3d�����j�R%��c���%yz^�j��Z�+�>��/����Z������(�qP�0)���h�����$���	9��\����ۀ�hYt��6�?���k�ɨ����n!/�O����s-���T.:e�ौL^��0��}\O˶*3��ofU%�Չ�S�q�xQ�n��'q#��۟*����ai����ԗ��1����k�#i�����]��>C��(e����8��i�}s��;�3����g���H�
���M%�ϣ�S:�=�Ya��
���%��7��e�=���0�7ʊ����;�M�@yj���ؗ�$:��G%O��"����$[si�)əY��T	�˚#%�?���Q�G~#��� aC������*�Ǯ�qt�D�*1Z�S6F�r��]s#I�ؾ7Q��x�&̹ȍ,�Έd��Q<���9z�Ȣ3��7?T�0�T4z�5�ʕ1��Aq ��zߤj-�傱y�u ��au�3P��H�JdW�\s����\P)�[XC�ࣖ.��+���nsx�.�:̟7"J��O=h��b�xD(��~[�>G�������Y���y^���)�'������g���� �0�Ul�NʚWs�������밁�WM<�I^�R5=�1wz�~ڡNւS�ā�A4���,�k�������9��H��(�	o`����3�8 Hy:Юy.��/�u�r���-k��y�QRb6���0]l��DT�y��۶+B���Ou��ƾT�h�-d!���)8�����D���A��^
o��!5����6{{Gx}&< �dq�����LCU7��<ؕ��<�����36���v.c��-�E6
`Q���e0!=!d�͈}r��rIco�<k%��P;�HOP�O7R����q⳨�<G)0Kc)<�y8�_z()���q��(��u�C(��+q��>�7�s]��<�8∤�<j���H��+^��4̏����vn	Ms�vUu֮G1�<��˱u��-).*��חU�0��c�!�)L*��#��q�� Ti=��h��<��kyP�*� �lTMn$>����.\�Y0s& in�jTv�8a���z����x���x�{�e�, Gw�M���_b���2ř��I
l.���0]1�n��"���,lI�c߉D&�2�yQ4����9�d�m�	`�]��#vM�H���'�ʚ�f�szM�t�t��r2�Ф0p�}Im(��j��i��"b�f�}&"tS�9����U��ɍ�8i��x8O+��!��d�	��GΗ��6����R��1�`�����/Ĳ���Z������f����H�Ɂ�KS>������*��eR:�3����|B�Io��4�w��k[_�h[�����֒&�tSFt��=�3���OK�0e��[�2�����ד@���0*����
����rδ���=����*U�<4x��׼�?�Y����o����a�{���}��/�E�KY�a<�@	N5\�z?�:Y��^WD3�ÉOdHt�t�&�K�z�"���Zy�w�~ʸw���f�:��[hȘ�Ą���#�=G�����(F^�w��ԍ]���A�8�zј��������<�Æ�}��J���7wSy��<�݃��x��[���9���Ҋ����WШ*��]bqA�U%ߩ:�����]��<�O�g�ެ݋� 2�1��j�Q�@ۤ�ՀӁ>�S�)��8��[�wJW�(�������o=���$G���#BOh
�Z\�&R,�>��2 vzۄ�(^��n&�o��(1svPG�v�]#��c�Q�i�v��GM����x