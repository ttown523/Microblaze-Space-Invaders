XlxV64EB    5d01    10d0�Z5Lo�X�]�dZY�A�TLCr�j1�<�u�rI:��p����9R��c��Ѐ�5$�L-%��&˔¬X��YM�	��f�NY���#*/��]�U+j]�GJ�^.6�]3 G�|�'��Rw�!=��*�����AJ�<�:�cG��~^�M���µ���l���0X�g��w�5���Y��,�?{Ҩ�_�2\1��Γ*����=8z$��U��G������З����j�9��(N�� )�N���ky��&�N�sۆڠ\� �2�&���(`���p���8�{�X,�ZYcV�|� �Bt��Uj��s����h{�V�-�Y�H6�$��<����;r�Gl�ڌ��8�Y៳0�ofNo汅3���lgݐ���o��	��PEp����JOA:�8KiF�� O��'��{����R�1�E��V��Uѕ�:Q��6ߖ^xe�/��C�nG��_91'�T�����,R� M��e8}g?~FQ��'L+[rf�$�yZ�}��L YN�Z|R�79�󎯧�^@Nn8(���s>x¥.�:������	��è-2���&�&r�GcK%��GG��%d�U��	���F<I�6Ц�+%���+lXݻј_���T�a�%6&j8���H��2�T5'ö�?ӎ(�҄�"��� �Oi*!U�����z-�2� d����0��F�	�3}�=�k�`S�p��f�?j7�>N��xE�]hl���F��P�T%�/e�y,�~Ƚ�$��]>�>�ZZ!��Db=�8��o<��.|��L2x��H� .��\�Ș��h��S1U���=$��-Ռ�Z$�1����|���)�T��g�/�˕d�q�%D�L�"�����|��K�SPmzj��Mp�G�;�5<ѓF��%L�9���E�ڜ]]Ʀf͖4�Yr�:]���kd��b�])��q=�RS%��X��(�����atI˫�}���R�n�a�Cy	�%Y4�{	�w&��VqvZ>GS̏�b{{�U:�����b�i�ϔ'�]ECO�ݣ�ݬV�q^7%�` �����{)��r�i�E��8�"{n�Q������^�d��ެ���"�`�H����+{=�,�ػ�U���Q�X|�{R��=C��T���hIы,j[>`�����̱�����h�}u)�`��q%ܯ?6��`:�4�7c����}��L�j����FlNÄYa��r;'a6),��Z�}My�ʯ7%Rŷ�$O�93�cN�C��j���zJ�,e��ˀ4S�t^V�8�W׎Z=;��<p��J|Ȱfۖ�^��� �]W�Я����Mj��G�A��Z�Bڭ�G����	���X(A��G�E'�S�D1kɃ��Gz��\�@��p���8��x
����	�����;ey�J]O�Ŕ�s/,%rPK�Zt��ż���kbٙ�uQ���Yأ/��J������ۮt�Rf=1n��#!ቅF����^`�ٞ	Ȕ�N_��2���y������tgE\���"J���Ͼ2�z�
B%-����[�In~��*��I��i�e�m؄�6x8`"FSg�y��������:�A�Ҧ*���:�w�j��	z���AX-��$����v�?I��i�bӭj���������@�B'S)�c������	��%�,�j�gr�L�J�	�ε=�f��g��0��4�i�ƫ������|�{즳������5��IA|K}�� )�_S��ҍ䋶]�.���� �� Ǵ���M�o�q~�xm��U��ݖ\6%���g�۟���v�9:�0�P̘�xC�o0orþ�y񱐚��mj��*��&1[}?ه�"j�`�i��PO�s�
rq�H�/c�ɢ�]���<z��i�\�+�s+;u�����.���0��M�hxS�x�3����|�����>�Q�����`�Ff��cj�!3��Hh�/��;b�U��4����T�<�qbz��8��^ĩ�YT�-[ޟ�`ɦDNc��X�+{-�	�OO��/�����p�.	�v�7DTn�� 3|�-��Nk��yqF6����s����$�Z�WQKP)A*��`X�N"���7>h@���{�u&z���
�W+�Zq�Q�^E�4%P4b��k��2�tJ�ߗ�j��_�=R��Z�[����UKm�c�3�R%��FR=�H@��$b���ꖃb�м��5f����$
n���2�r82���� ���J6�d�����,��Q~r0�JM�#v�%+�����͆n��"a������)U���i�[s>���RCL1�(6Q��_@{��DЪ��n(���� Ac���"��N{|<o���wd<��t��>��֭.�����j���|�a�$H�����Ｍ���H,� ���k�}�`TE�� Qj���C_zku��G��XJ�F�к������CP|���gN	%i�U,� *7I��O\@u�Z�$`��:�����������m؁��!�~lNdʐlԃ���X:ۧF�oP��.��r��Gkш�������}�,����YA卶n=�.��e���zd89ȕ���L�~9+��R�6./^���y�8Y$&9��	��Ze��]�S�ބo	U�dMy�w��&��
�9�;Et�^�}@����
򔱺�u�JF����x$�n0�����NY-��/�緶�G��eWӱD{~�*�a�c�F��6��$����W���Ϯ&8��rW�F�㽚 �f=�*��7d2k��^:'d��и])�&Z�z�_-���5r6 �OHs� 
����#ʎR��L�zN�u�a�l"d_�pOG�tS����>��	uF��&P�)h�:;���� ��qŜ
)��a���k�id�J����������r�Ԡ�T��qTb����oF���^O���_c����&1��L�d�zī�/+M;��弢x�F���AT�L���E�-պi@��kZ���y�وʝ��B4q���8׫��D���m<�}C��ủ<�-�=���sy����9Z�tw�TZL�{8A���Y[΋F"�*�8<r�\ᤞ:�1��+���A��}�V���et�U�2|��4�mi ��������0�B��K	>��S�_�	� ^�z%����Q�~���G�o�v�uBi��318��Qw$������듁����'I`�|��>�	*����B�����j����D�>�����<~���3�Rߏ����&���ڥ3n�L@��Rw�-���?���ʀ6�P��ϊ��z�R��r���%#�@�x{aM�����c-3�������S=l$~��K\�f��@�߬%c��(I�S0�����S��G��id���'M^�e5\%�t�K��v�*q"!]���;�MZ�>n'�jO&���N芓���ȞSWh��j���q �R�"�~���/x��IrSE��u��)K��4�|��k{�0�� �0�n�L�vȽKu�h��܈�pSҾO���J��>''47�U���xX�c����-�S{Jh����J /nAJЀ�1�'�ľ0��������@�`x{�9��3t��m�7$��@����b�t��
z�Q�����7}�B��
̜@:�c��3ŌO�����6�Q��dA0��:z.����Y�1­��n0�\>%���N#Ӟ���qW����J�=�-X)���e�落�|�:@[O5<���T�n��h��"!+��:rBA�|5�y�Kf��>\w��V
���3���+J��5�Es�@�%z86�n�n������Dצ#�PEպ"%�=5=.Y����B�+�n������}���x�.̛��v�ٳ�W�R�o���K���8&):��f[c��aqɂ�q�r��IT�i��3;����i/O�*cu"�T7f��~N\S�D �s�����S��\R�������|��cb����N��,W1UH6��":A,���V�z��X�/S�[f�X竆�ZR'���0*�;�*2ꫴ� @�l^�+�??D�c�h�)�-/*��#TT��;n����_�B����^f�2�a-S>�tߢ���#��! ��NkvҖa���jzl�㟊��~*:D���F��l�mHxF���!U��C�8B�ϟ�J���~�!�N�?�,m�{�al���(UU��tP�O��'.3���.��OW�Q��J�)Y�W�U�)[XvD�