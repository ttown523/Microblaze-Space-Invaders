XlxV64EB    1edc     aa0#h�Ԋhގ�.�x���"	M���/��>Wao^�B�$�a\z�_bO)z����ҘF�D������Չ������>��e�@$�t��kB���A{_:�q���M&��ph���.� .�M���QB�G�W.��9P���8 �w:1�V�pyc{~%�������fg�B��5���m-��$0���%v��|k��Ky�@�Ǫ�T
Ł�z�]��:�H_ �,+4�<�a�?>!���YL�4{UJ*�̨�������v�U��b	PӘ�U@��9�� b9p��,a)�{���Ge4uLh}���`���2pG륐�Z̈��mQ�Ck7lΩ��#�����=u�-9W�jxmt ��H��کL�y!�p#`���܋p"��,�q�#W������4���d����_�o	���/血��DL��l=��_S�y���1�H0~�4�>H��7��b�E���'.�f�X2b!a��e�����w}��0��TVL�Yl�߫$���wB�hvϩ�O&�(�O$c�8�^׏�i����>�#��1�0�B�+Cp�֗�iZ3�_�5�c	ӊ�����M���L�"�^�.��+@߅4O8�0ᒨ��/l�W�D7�F��#G���#�K���,O�3�Յ��ͥ�=i��|Cs�*�w�i�#�&�n.��$ʅB�Ϥ���~!{sMı��Uk�S ;�I����������n/兆H^���	Q��2��X��&L����i��O��)+��z|Uc�A���BSOs��� Tg�I(U�QhCQ�����L�[(ܣc\,�0qh��K��/c����t��_(y� B���Rg��Z�/��*"��@��ޕ�Ɠ���uJ&ѩ6׊]��w��o�/be�����'.t.�O;�������i�A3��lY�1�@�9N�;ފ�G��r���Y�v^߀eMHd�e����Jf�`Ԕ�����qnD���2��rՁ�˨���u(�p��]WP��U*�B�a�P��7�C�."/\W����{�Kj��f;9��c�8�n����a���w��.�7H�F�l}3s��J�T�l�pb�A$��l�A8F|E�U�"=.;b�䴜i��B��u�&���6��u�� �~(��Ԓ'�eMH�2M�ڨe�V◓�I
"o_�4��L�.n:z�,�KҀ�Mo�蔧Z��Q��FIUڅ"�ZF�D"��ʴԊ���>Ă��x����7"_ʰ�aϗ�*�$=2�/U�,9�Tj�6�,��Խ� H>�8��C9�����+�`�^w����Y�.P�X�����aӨ�1��TX$�mFK(����W�|��<)C0�u�a Zٚ�21�o�Âa��G>>�iz�oK�V3��5#cI���J����U����/��k^(��}�jK��ٖy���X���A{������ \�V9�j�N�s
$�Z�t.��*�����-�Ȗ:T��&Up�c� [dC�1١]��6�-��}Y��Y�T�������{�����\��
��p�ګ���%�lMs�R`�X�����	�z�uW`�MB�����(X=gj�i�f�*"�����3ϋn-���Z�&��I*v!�v��qUP�cx9�r��-���hHg�����as.��laSא��-��/Y�������a�����pR>���r�H��{S��ӌ!)��.m@T������R��7=hwO)��'V/C�;���í�	B��dG��á��R:*�:��
w|9ő�e"��_7U5��N�)b����t��:�����+����.�����E��kVu�o�v�|���@�����_e:���#��sb'G��gEnq�׈�0�a<��mH�E;f����ҝ��B�]ީ��ua����*,;�F�_�#��`�^]̻g�k�Y�?Â��A�}�Ǭ;���S�a&7nji�1�$y�(�Q�J�b�9�d��)O�K�/� � շ����O��v��ܣdo�)���#{��!h��H,䒰�}�y��G�Ch�c1z�~iyi��0Tn��+8Fh�"�&��-y�0G'��q������V���h�A� �|?D��<�Ʌ��$��T�٩
צ�%�
p�o���SΦ�׍��j�2��琼���:�*�$���ct3S���]n>�H��[N���36a֖gƠ i}���2�����C��Mӊ���w�#|ȱ\zv<�b���g��/O�H>۲��'�A�J�!Z�Z�<��q�=/[���8�m��(���0e����Ei1Z<�d�Zif�݄�������p:՚?��h�Q���6O�y���	۰�K�
�Zh���%��	u�㫵${��}������P�b�"�(\�eU��)�ݸ���o�O���]8����ǀJ��nY����W@1��� ��Qu9}�	�f3�c[���sLA�X*���GPB)Z�V��~���	U8�^��i��Åv~��q�k��C�r�O䴤�)�7����ZX�g�*�:�����2��V�d�����B��x^Dn��c���V�������b5}����^�b�f* �"h��ƶO�Jяk7EР����HJ���ʯ3��y���g˚�����4&m���ű�n���C�5;4����U���.|�=J�H/'�*���K頼����rܫ�k��Kr�