XlxV64EB    3a3a     ff0�i	,�2��[t쪓y�:�g�q�T�s\Ol��P՗��9�,�b���<[��Q~ʱܷ0�f���N(..�n`E )l;HmYO�����T׵�ɏ�����(�n1.{B�@t���~i�!{����o�:V����9�����)%�	V�%��~`~����d�p���b#� ��C�-20�t��� W�F��w��}P~�x�P"l��)�|K]�����g�e��2˕�R��i�D��%ZZ��.B�e;�����������O��2x�&�fi��$I���e0�_E���x F^���&�zd=WѶy<"	��'W��|v���03�ԭ+=C �����b�L��h�؇�4<N
"<Ro���aй|wE��˻����$�'�;J
qZ~��=� �t�Vu�c�f����b(���8�ǰ:�H�<��'��������e���k�!���-̦��i�L��#GV
��ކ�cؔOZo�%=��~�JF�(F7F�,FK���ǀj�^X/Yg��I�N�i�[.��s�0#7��=��a=x�tVƙT��>���rO��##;�̭�AD�*���Έr7�{�LL.�4�6��_��%������~L�0�Xd˓,�-��ƚ�w-�pN�����G;����l���.&%��ja�����E�+E�N�F�<E����L1��c��6|R,�
Om���ds�r�G���l�� �:�W����jv.�gj�3��&u1E��=qт�'��i�w7�����_8��$�A����1�`"I�3Z�"��'b	g�h(1��zI��n}h�ue*S�A2�sU⧐u��%9��l@<�@yo�C��u�VA�'��s!FP+�_1��X#C�~v�o�
r�leTA����8�>�-�6#fwK^��}0��\��Y�(::8O�Ж'si5Uq��a�,�Fv=~��E
��8 �;]����d�l*m�/�L��9�"9�r���^[
_74�Rz�R���S����z3�~Sz*��+��P����B-���T���	�2�`#pNX�w˰S�����s����'@|�7�Y,f��y|��q8r��
�D�\�����|�Xl�{,eA	�blO�#�fݵB7�!*>��-q�#ꨛ^�@��W˗��K�7����c���aXv?��TN�.?�q�Cߑ��V�6\�W�y?����羻�Y�n9�]ծW��hj� ��� �]�(��������/�Ш���R�!�-��T �3]��y�#.*�ɖ���7�sy���[��b�B�IZ8.�=d��ǰ� I�%��N�-G�]������^�$k�uQ^�i	��a�w�N�3�-ӷ��݆׍�|�AYe�D��M�{M�o�-t*�����fyl�ˁ���A�?�K�vBe� ;ԟ�G�,�F�K'hζ�RV��F1
f��+�t�UfDx;�6��.s��p��Se��c�~��"�-D�-(����C+h�X��J�� �/բ"(*�$��f=�%	��pq���.`��տ^�fF�Fi8�֦p8tOm������>X���i�<yc"A�/��eD�_^U�fQ�-|Y�AWc�G�}�u����qsA!��+�_�Vū;	[1��S��r��Mx>�qn������*�L������͸���yߏ�b��yR��
�Xջ�΀�W�H���M� ��k��Oc��X�|1i�\]�B;�mVߪ� �Čj� v��EwT`]q�y��"?��R!��Z���9|��_��f�d�r�٪� ̉kl
W�s2zG�B
�X�N�.Y� Z�����?(�o_��H�n���	 �1,�V'�����́ų%I�m�Eu�ϙ{۱��0{���0\�HV����K�<���R���Î9�����(\a#4Gbq꜍͉/��~�y ���@ �(���9_E�n�4�;��s `i݄Z���KK�à���}�KA_�A�v�R�(��W�*oń����b������1�ģ��81�{�p�biBU�]:���q���|`�];KsC^o��yc��?P��o�i���-�kMN�rEt8<F��΂������i��e�ITH�Xn]���4{8Vr��6z([��k;��C��,��e�:[L��?.�%�{?ʬK0��.1���&W�F.�ڒO�M	�v-:���1P)����;Tج	�:�mNt#�-㧂q��'̮�k�J4v�~qw�����26/�ҭ�9�����(��6�b򥶩���i��1'�f��a�Fu�n��x~�賃BV�JyW�RT�]���&���Np8���:�v!��!����.��]�`��N�DRu����O���f���\�a��h�8k��	�A�Z3CҽÂ��<)��0��7	Rx��,L�T�p?�d��a��Oӎ.1[��ӗ��;����RP ��1"}X��|�bφ��� �܁��2�����'ڱ�:D�e�`�`P�k]��2S��*�8����߹�F���	1�y$�a~�������F�m�OC.l�d���`!�����&���w� 	�]�)�[/a�p��9�4�1l	o�d�֍\jO��|_	� d�,^�'?Q�/�O	{`�&�x��~�?YjSi	�q�N���"펯�M�L���̥���_�E�7T�v�7z�U��+�Z.:�v���Sr�b; |�:!����̢���[ծ�0�h�O�iq`�P�0�Pz)ld��傇p���rv�=������P#�l(�>�hN�Jd#ู�B��ul���EU���&2N,?��%K�_8�����VM���3�
��S>p\</��뻓z_*�����u���d�NN{�q�;`����9���+Z��4;�5Y��
�P=�9�V��Ca��uf�#�-S�a�V+�TE*�c[n�&+�
MC�Z�^5�$e=�ON(k�oo	�Ϫ$e\�i(.�#v.C���/�(��	�;��]�>Vٍ������3�0�2��KAW+y�ڃFD"t^4��� ���xy�X���h.mw�w�Xo��[���s7�����UM�5���'Z8`�}� ����2��`��]��~�̓<��vuW5��%`m�u�P�4�`C	��������Do,,@�����)�lj�9Q��f|�Y�����#!��S3?h�hћ���=ǽ���F[���_��:8��RגJ�H���詊����56/SIN4�6���|0ykF���y��v��+cv/�O�=
����ci!/O��m$��ʝ�Y�� ��*���~�ΐ�AL�����J��%	���v���QL_�	>���dK���G{��X�9�5��-�랽>�C�S����ia��gRY�l�U�=n/�3�}����ۛ�d�B!�Yk�V�a��$��q�W�?��32���7&�A\Ǝ�hfc�2U�+L��4�ْ���=����Bq1D72%���4�\� �)ռ�ͮf��y���O���3g:cl�a1���JrS-*xbPX���I_�Ǜ"�t°��!���D�R>�cYw���B���s:c��=C4��Ƚ^u��ã3�t���#=)��S����a.�j���S�u���)�n�|<B#֗�}:�MN�i��&� ��:J�u[le�bFVe��O������e:ʼ�|�X�7�"�hY���q��G{w�-�iPh��N��M7�f.X��T���k� ͨ����y��2�>��?�%S4L���|)Fcr�*ZF}\�O�=b�T��p�5ޤ��>��J��
��nh�nR�ǖa��z�d3w��O9%�t��AnQQ5�l���k�I!B���Z4�F����۶�f���V�1d��s�	���7�WQ�>�Jr�D?�x�;!��k³��5T�@�j�)ֲ+=�Pl�P	�t`�!��K��g;6(����ER߯���\�v��}ĐX0c���ׄ� �>)ϭ.�T~��@82�T��,����W2x�_hɶ������i�x