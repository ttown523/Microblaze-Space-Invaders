XlxV64EB    fa00    2f90T&����u)�mk�9���o2�v���l��,�M3�7���U�t���;o��ڌ�g�b��Q�_�i�f���Xe��-���,�E/k�o7�q�g8p���3>�i+J!D�������1�"Ef��*A)�Wx�p�n��kҐ��A8Wp�˭�A�P١�f�I`f)�\�u�u��_��[7��w���}�+��$L�(����z1<.fA�X��Ʀ��tT�Z��@]P����(�8�QD�c��1�f
��)#�NKz���/�l�hg_�������2g�x���71r��}�c���:#��k(M��_��VY���8�$$�8����Hc�J�4��Vi�QY��(>9�2����kN�o|��S雑�]��0�,������T[��E~���EMZ�O�ت+C"����b�wf��Y�ˎ$��p��a���I*B�D��ݢP)?[������~��Nrk�e�jWw��Ƽ9�+E*=�a`~5n�M�H�����P� 4B.iڴ�?ĥd�#���j�<�������s�����w��}:vwBHA�+1�"f�%�S���e�փ�ۧ�f0�B�X�6Eo����j�Dg��*.��T�u��C9�p�#��d� m��n�¡^����@'��U�<��7�\��\���B��I�(9�Gg!3�H��%�=결�ܟ����c��N���m'U���X��ZPlX&rR��R�Xh��ߩDY�e�l�?_��ґ���^w �W��ƆdJ�*��w6ز���lH�d��	�Q@
��2���n�}�����|�	�}^��=�"�|�l�V;M=]Z��?����HH8�&�wJ\���o�j1%�c�]��)��)D�{o�Q�5��o������aI����xQ(i�t�iv� �E��:����,ri�Κ(b�A�9�i��m�J�γ@ ���Isp_%��K�z.�t˙�K9�A��n3����GD�
f�,,�M�L/uj3�� �Ы��� C/	"v��%흵�{oT�ΟT;W�W^w �p���O��Q���3iL��*����dXi[=Ӿ�ȕW��@���&ݮw��;N���e]}�hV3�`�I����[��n��]�/�A� �*ͤ�j�uUI�7�aD����j�&�Ǧ���&a?:�c��8��A�z�niX�|��>���s")f(��O�"�>ֆI���5���K�7lhHը(ֹaG�����[=989PՖ�9���o^`��������rs���ˬBk�((��H�A©�To�+��(�����Ck��JPB�aq�a�t�3~�k���3�F2���*a�����6����Ѩ�B��t������IRNB��@�ꈷW)W����a/,�}m��U����c���$���:퓈���A�h������㜚����F1��$��mw,�)/yk��u/X�bs���UG��7k������*�̱[伌�����֠��l�}�G��W���M,�j|L4�:4O1:�N�P���f�q����(ɤr�PTz'���{b� .�A=�o�H�:�׽�䛙�M5{K��ԮÃ\ @��.K�w]4��6�H!J��[�76v��*%�4|�J�j��f����2�����_9#�Q�^_
��W�B�ɘ�z�]5������l<�nȡ���H��#��~�\�{��0{�b���b����������lŦ)�UyvTw�ʵ�)h�TeO�������B��]1 ĩ�\��лQ�����i�6ޯ�ЎZ��y���{�����������Q�m�7��l��Q��k�5�6ܙ����1�q�n�Ť�?�k�B;C���}O�J:���*[�]dQ��8�ѻ<�|�GhV����B���+RdvBX�c��T�B��?��G����CFff ���.�nGJ���d�6�~U��j:\�v�uL7L$2�[YnK\�rpnP�K18�!�r
(I(ks�����kRf~'��b�f�13��-��r.KCD�ȅ.' ���.m�^�����7%B�X $��Y�e��^���n$������05[`2[���{�������ԁ��;"����Lz�k�S;�Wp��ء@S�b[ ^J^l�NpS]�	��Ϙ�	�����(�C�Uï�k!��k�č��h�P�Κ�Qc)��t�h0���^_D$A;M�0�}�o+���~��p�s\�����((�yp�A3�����S� }z�cH�&�z��z��~O_2/�p�#��	��y����{�`���wd����v�0&���LI������;\4>�S��_�$1<�(�_�x��n�[�	0aZT�ι�K���s�wbFh:#�䤴3yC����n��W�Kkw�M.Sa[�]�-�O��pN��>�����&w�ã���Y���!���U�P� �O߂,���,ֺϵU}��0���RQ� �[��k0狯6!g5� ��C)̓_�`d��		�C���Ӕt����Id=ŷ˫�B.��L���K���Y Y��kn��\E��dK���H�J��,�/^�W���o;/L���ɔ��Ɛ(3�>_�^�H"t~�������u_���/�⌞;i.`���STl����TW����W���xFub����x>�7�1��^��"�~w�ח&xa����@|�,�yH���_m� ��P��Um�������ߧ'נ�9�(�����0��Y�i�*����}u��FJYڈS�"�t�<�����W�E��@"�يcEр�Kv�%
n�持3/�O��"f�
�T����>��/0�Q~����f?=0����J�7��25��)#�Z�!S�`ͅ7o�I)gR����[Tu^U�ѹ��X`�q=Q�"��� �\�EWI�(r��Od]馿����V|`7�{�g9}C�={U)P�������q�~�U��y�s��u_���Ȟ	l����K����`�
����跮s����&�ܿ�L�C�C�MP���Q����F�N�e���}{x�O&?���}������Jh��X���:�� ��Q-������y���7Y 9����u���70U2"ƹ���9����u,6Aͮ���YsTo�YD�H^��jA�� G�=�q������7s9�0�pA@���+�]���~2���1,�ю�g`7\��Q�l 9�/�+.����Q����N��Y�����W(�i��~�"cر>hP�
IY��c{�����ݏ���|
7P{�|8 �e:��q�{�73�྅��y�]A�0kC-��2ԜYѹ��V����Q���1��	^y��|0����.I�dAD��pV�٧�	��R c�
k���k��V�~K���x`݊O�g]�
 :���Z1�s�]T�7��z�|�������<�Z� �?��,�5�(�RW�;Ǐ�*�ɐ�ߺ?[��ȥ<O�tW�+vQL�x��kґE��޸�i/	�z
˃�7�ʅ6Q��D�{Fn�`�u�$ ���ћ5~��(��Csj��<�|��ђo��V�!�ajv�AG�rB����y;�ߨ�ȩ?I
1]v�D�=Z(���X��e�!A�;�;*���'��!�����7n�CD�}����ma���c��ٺ�f*������Y�$A�8yHU陽[S�ߠ�4m;
�Qw�ؿ��	Ƙ�v�A�t�Y�\7(�� ���Rm9�߆-$]#�������r����e�Z	�0�����½��vVyod������,@��mAo�T�tI�e�v�}�g�zi���ֳC�I]�q='�˧�J3��8镅�"��Ʃ{�	����#��dJB�<�*��5Nz݉���Q�lp�`��=J5�ٟ���,����/��%u�H��U�(Ov?�q"}�kD�Z�X�^�<����x�k:%��>t���o��"�Đ�r��{��d��	VB���NF�ԩI��g��O۶�Z {
���� ��pK�K��ޭ0[4@�O���j�V��Ʋ �q�S
�Y6((�jK8�x��I#kEK�*iD� Y���"���]���S�tg� aеV�'`�H��f�]g�R&�?�{_�H��)�h�	`���j��|U��o�¢�ۘ���F��+�!dw�~����e�A�h>�yÿ(H���XyxlZ�SU�)I����ȇ&^�J���qt�V�����'u@�����`
�]jd�2�ga'�j�}�[�����5<|�Kk����au��(9h�fxVy�
�"'�����J��eU�R-Z8]�ρ���5uk�r�&ݤ(_��������b��Zt�g^���ȥ��a ��p�p�����l��n��-/�V���웕i��غ�g1����_cٙ�5�bؤO�\��b���T�Pv[ƾ��u��{o9�&)�?mև,��շy��D�W�sw�tp������R�MW�qt%���LG����>�<��J츥Up��`��vw��.��P'c�p���G%�Q�0sR�_0}�&ED��g@cy��:���6p\��:~\�>{%�����Nԯ�~�p�S��	E��%9;��S���y�)��'Ђ�ˇU�<ߒ#��}"��2ē���sF�6��2g�3��kK,dl��hХ�my�~G���?.�6F_롅����/̨�)�9����-r�q��"��;pW����eP��t�	�B����$�v=��"d��}Y��`�A(\�׏�Jxc����N�bP��
;?��\�',QB�}�}���,�n�����bF���:�E�!`��O��߻�ޖ4�U����	WB`풖���ʮ�����\���!i(�`Rp��E�)���}yj
�������L)ʦ�� �}�A�S0@.�N�n����+�Mi��r�Q��񏠾{Z@چ�DMOO�����b����1Q�Ru�Jf�8�J��Ix���d
�H��mv�][�`���b@jɾJh[�v	�*�r�h����� bĈ���͞�4-����<���f-�G��Q�'�zMMW��ߙ~��7��'WeH*�F.�����Hh�����Uü>ҎN!�c������Գ�����X���d�(JDR�A��ĩ��&��\�3�^�w&�^8��W�x�G����HT��:�g�ϡj��/�� �Q" � (ft�S?��}��CU���1|�qC��ΘDR�6*�=�׾Ӣ�\i�g��I;u{7�~!�,��Y�5F��OW��op��-�'���K��mUĆq@a_u:�����CNx;�)�C�ܰ��(���O��������x2fC$�@0+����\J�@:S0O?��CcLm�xQ�>Ƈ��L~~�kdh�Ci�N�[#Oܿt`a�(��}<�"����y�E��tl�ҵ.L����p������;�� gI+*���b���=/p�<�����3|!�����dC��hJ>�h�d���Z�}��bCW��_q��}�����ryPg�o���cb0�C�0Z5iykI�rቸ-�7ͧg�Õs��H%u�=n��x�Ne>ר��k�����a$�u�֪$�18�'�V�E*(�b��sM[ֶ�I�'�B8�Ka������n�]������[r���V�9&���1?6�O�uf9KM.qG��r	W�@t���*�d>/7��Ǿw�?ԕ$�|R,��|��������m����e��Jr%%ͺ~X51�Df�H��Xj���������H�r�l/�|=�Z��������A��j��p�B�́b���#׮�DZ�~�N�暑���,�I�R����R�w��{�V�Yҧ�m�T��A��(�Zp�t�ȧG^����VP=Z�����j}Ǝ7�6/�]A
���R���Rc�)_	(�.	�`;G+�|����fk6�����M,^$ӣ�9TX��m�'�Sj���2ZC���к�_�2���:c�#�ȣ�ցW���w�@��{ �3��9�x��$�h8{Q%�]}�L�͏��3�&�f�>,)����3�]�I�'����:����e�]iӖB2�o�;�7�������U��?d�J��K#:tߙ�+�¼z�=���A��M��7K���z��;����?6C$��G��zf�~���,�0�R$��)���v�������"*���k��b)�1�E?�)cl�^�=՘��YmP�mM�f��d��jS��wo��У;���d~K<Mž.Ĭe%��7�����0�ٱ ����~b�P�z{��>��a��WVېGLݎ��ШQ�m��%
��z�⍞q�=���,���N>��?�*8G�c8d�����9� �����I�5M,u2REh��d�-�����xX���M��,����^]\	-�v1"�4Пp�$a���('m!�W��N�3��Y*�	�F5e}�&�?��j�Wbv����sRg�p3I��xʈ�Y�zg*�3,�rѰT�� �z���v�h,�6";�aа�eX�6�Nf��c�a{�\����8��ҋ�7Ie��y�E��p���F&
�NUe7��)������u�]���p�3Xk' ��gS�gM*���u�/Ս�.��|p���n��#�ڝ��XD#n�X0u��y]_W�]#u���ׄ7N��׼s�r�ǧ�sIt��NcAݏ�����b�S�mo��,�$V�6��e{m�j���.�����qe�Ņ"�k5W���pzB�zt�B� 3λW��/�yp�3:��
�.���F3M�	 ��XG�Y>��������e�������-E�g��N0����8��d���9��G,��.v���7ǝ-�(��`��ڦ ���Q� :Ҵȯ������
R��$�HP��q�N�>��'`�E6-R�!*O\��6�7x��)� )�<�OG�z?80S��D����Y�(���5\,�?t��"
P%Su��y��b;�7�$�*�5���2Wk��?�܌6䕀�C6'J�O���I�5P��h�T`�
`b�3��!���������/9�������
��t,�j�x��k�1�U�M6zb���V�]ד������~��D�Y6;5[A�j��� ��l�h0�@ܖ˲�0U2C��:��w�M�q���4j�#7T&�c�Ԁ�m`84�V��KT����	I9���?��������8��>]����d��6�5�jׂk*@2UI���B�f��W겧E�Z��<$8�XjԜ�$T,~�y�� �4u�����/C۟*���y���߱��*�����de{���������ʅ� ~d$iG#}R3"<"{��HW�k��Pp�~!^�aɟ�^��L���|����0� ,H�e0��!^�O�%(C���_�Ւ��u�>���l��0��-�V�v��dS��H�~~?. JK_��\z8֢t����z�����O��J�x�% �@��F�(&z{�Ja�f�9U�O�rr���y_U�{���ՌtO�<sF_�+��.����|�p�%p��+p�0�^���Λ�b�_YE�5��OyfjH�+�E+� o7���|���(��Ί�F����J��|u�Yv�1�7��PA�&�@K�nƀM�%y���ñ0x���[Jw����E6��`4�fp��Ti�F� k�0���llf�Z�\��uk� ���V��&��T����C0j��5��7k����O��z��Mm�<|NG�=�JG���q�c�s��$�]n��Z��m��8��n�\Q����8>�V����It7���%L8�.^�ਤ�E�� -��w�Z��?��[��8GUj��<>P���hNƷԌ{��j���iz���*V9��e��&�(����JM��ӏ�>�Jv�c��HܓR�]d; vj�~�����n��}�77tm��ն�F�J���`���h�;&3����i"���`[�P���N��a���Li ss$����O�G_����܀M�G�L�?2P����k!��ҏ`�dƣ1n��e�,5�ƍ'��/h +����f�q�O$� I�i����K�X������!/w��z�\�P<�;V��*5��P��V`>�2�Ep#���v�e��B��*.�#XϦ�����EG���?�	�B�s��3����/w���O�pW��	���~�%C��-bB�����6�8X�%�ﯻoxƐ��)m)��i����!:A{��J�^��L��~�E�.W0v;�`%���|Yg�}���M��:X��4�(橾�V�|D�x��L W3�t�-���e�ㆌ!o�zd>��aFH(|�[�~D@]i�w�8=�_6�#�_lW���e�+k�)�u��R�l��?RA���
�eT�
�R�w��j.���k�yK�F{���C���ә��:1b��/�Q��oF��-Mb���=��T��d��B��ҏ�W�������`:o��>�(i7�FB�o?C�ϔ��I"RsQ��=���m�.b����ms�rV�_ʿm��+�չEV_9�5��vV0�����PP>����:á���aD"a6�(��h�+��\�����"w��r�����+�?r�zZo���<2Wow�*����� ���P�!��8�_���r�|��0x���h�ā\o��Ճ����G��� "�����Q�mr���4x��������aC�/e1�Q_s5p�_�Ҭ��5Ȅ(��Ub�mH]h;rM~�T�L>Ӧ`�<�C�|9C�Kᢌ����b�0�D	��Ĵ�/,>E1���1u?
����pMڇW�*?H��Ͼ��-4t@�m�c�ѩ9P�����>�ieհ"��B�I#8��z�Q��N���Tis�OR�oQ�ݪ��
Q�Rs�$u;;�V���{P�:����&\�l��aD�W]<S6�C�j��5����?߾�'=�np��3�=�qHA���2��:P]΁��J{������J�e�I�!/�U��C!�Mt��O�:x�J��u<���Km�j��V~�}$�)*�4	'�e���h@��Nٯh���b�����Pg�ο�	Eb�!�>f��������<�?��4_�f��&8�2�#:��3�)x�>=�m;��>o���wEt�V�j	�gx�֟��ۦʒ���ʑS'|�7�"I�'�t��5�;�y�S/Up��ͮ,�f5c�����(~g�7BM�2�,Ѿ(��,A����RO����kP9��!�HZ�x���R�;�>$F��:�KR�j��}d�p3� I	L�P����ѥf+ټ�|{.4��Ւ
��
��8۷�!�����KQ�7�������p��+蔁�1���iw9�U*0���Ӏ$䄢��ѹ���X4 S�)&Hh'�����i$�g:�S����6o|�M,�������h{�����]� �(�kĵ{B�YM��X�ln�13���r�/S>T0p{A���*�#��Ֆнu�����l r��ذR���nZ�C��1M�ɤ�s���;C	2U��Q8�K����j�k�ֆ��������NPpΑ(V��=�m�ɬِ)�xg�*���s%*`)S�)L�J���B4�Y�/�ո���ű�S�S��G'�<�")ްA���]�ME�����c���#�	7�g ������n��y�H��3%/T�p 	��Q|IxᲾ4Z�)����	�iG�;Iǲ��W�T�s��M. ��C�''�7F�ZN�CU4j�gp�=1�8,w�zt�'Ҵ:��vG-�m�x���K�W
�n����W��A��,@��|ņ}!D�YN�P�� �Ά���d�/̜nO�r��<&7��b��u��?��Uh���XnS�I�C��d�����?�._���u�ʛ�y��.�"2H�!�^z��������귖�F⽡,=�)!f>a	�o'�o?�g���Dp��ѡn�u�b��#0743���#RL�u^1O(���1;F�:a��=��.���Z��8N�
�� C�IG[T��$W��"8�ׯ[��d^�"f��V�$��#ǄW$��c�чL־��z�t�W!Yj�? C�Ѩ)0Q� ��T�	ӹ�U��}.���cH7�:�̢�U�!�$-�����L�=�$G����9\c�i��+�j��#o9��ȔY�P%�H�E�	U.�Ϗ2j�<<QG~4 %^���r���m�l�wC~5R��Q�Ϳz����[��Ⳣ�+#��fK�.ҟ|�����_�Ӽ��}��s�,�u �t��7μ�b���_��%* �g0� �
Q�#:�+��������!v���9RO�?�e�l���Nj�z�\���/�ό|j�L�C�u�&���%l��@�k�r�裁 �C�;��K&� 8�6�n�;��"�h�^S�An�eqcN��d�"�@�
Y�x9���+�.�����g*�ȳ3}8�2�d�3�'oX#����a�B['�����R�ͤ9/�,����o���V�7���9��q�h�5�<���@S��R\m�앁� $��E
Y��CF�ЁɎ���|�&�E��RB�+�>ֵk }FA�a|��EO5n�0Ka�i�bQĳ:��	��#Lr����B�=z%�t���U��ϻ{�֭�vZp�w�GwR��wl��
BΙ�jO꒱�F�6P�����E�'7|z��4v���Aމm�W���]e�;P"Sn�����@8(B<0�Y`G���3l3Y��w������r����q����~OH�cvN��Ē�C�g+��K���Ƕ� ��f�7"������$��i����mY}��	c͵Q}6�l��N��<@�MS�#x���@��B��a�0ܓ~Iw{��GI7�"߀����e >�r�֯������������	~���ve�Z�SYy[�LX�� hd�G�s�|��9�ҽim�V�I�m�\����pbM�e�����𕗵�r��V�
ٚ��	�\u��,��������'Զ��ș&�u�,,��M�q{�v{�R.�:,�"u�Œe7�������n0� �m����S`dm%�'�ۍ���s�`S]XucwQi}[~Ze;����M?j)m^��'b8eň�(=䎪܀A���Z$���ߜK��*�s��m�F�􂙞]�/7E�t�@�#��%Ρwe��"����$~Ζ�T+9yd'�RU)m��̘6he��l6�0��:&n ����r87e�Yf����7:��%/��0r���C���ؒpe);�N����!>�e�҃�f39C�
3_�, ����'�~}*��-�ݜ�޸{Q��0~(�g#��|Ҷ�<?��ʢ&�H�.~Dh�p�|��t$��Av��}!��1���p��&8Y}�5F���]m���#q����Q�(?=��Di���&�0A��	ڈh �;_ř��� �)���!f*�;�M�,�Βm��疆:+�&3��/�$T�"�9!Y��%��I��ǞC̟PI���Y~�����th��w�ږXe���##A���πx�i�1E�QE�gQ��Vz5UD���t�4h�9h�Nwft�X��Q��-?�r�ґ�i9��J��<D����|� ��ϣU���QR롶��?�N�:r~�@�Fo�D`�:��Ͽ�ߺ�b!ş�00���S(��^�*������ƱS�®I	��bd�����Z0��;A�(�����Qn��ȓR&�^���Lk�z��4S�6�T���s*��q]IN/�t�gnLn=y�Em���q�ȭa���D��G�j���!HQ�j�]��V�K�6cUEL�./_�f�[d0���K[!�TQ�����/�`��X�D�?�/_u�Xn�����,b�}�Q|���7��fT��(�c�#j@csg��'#c�^�8��z���cV���E�Y��q�o�Gp���ƈ(���iw"O.�@?ѥfF�ҙ�x
y��sbYf�pba�
�����*V\�';��;��A�a�5v�ѾXlxV64EB    72d8    17d0;D�n��"�����)������~��J|Ɠ�[[�"�Y����2�ۉ�B5�����o�2���,���M�;���T�,.��9y�	gX�f���5d�3F/��v��$�K�ua�uIU�oR3B.���,>���"����C#}cql�'�^��ڠp�G�P!L(�&Xz���:�y02:[4a������jt���Ѝ%�	�����ܰn���&���w���(�(�n�䈻4�:����ܶ���~�Q���8$ Z^��.�~}���MO��]�%�������[�f6��^�:�-	�/�����(<�6�~�)���.���R��dn8����p����j��]�T���j��zc5��r@y���硾�^Ly�����n���H���|�C�@�����S��a	)��.b��x�2����=v�h7�����EMH޻�c�-��4J�!�ԫ�I��Ɔa�qC��9ڛ)AR���cC
;�k��&w`1��L�>����ϤPl���+�݃y��C4���I��P]ڷC�p(���̄��O!�2��	z���i��.����ED%����dބ3��T�����c�H@gi��)��?��:ڊ�i㤿5vD�P�*�ޖd�{BߵT,�*5gl$�M���=�D1��q����g��F����i5���t?��c�(0��{Ek������$�(�jH����`��?�j���,}��e��C��8YT�ĝ~^��T��LZ|��ł�k�8F���x��P	��ȥ�l��}{��o<��x��P���ѲTT|4z�9�`�����1�E��a�H��M�^�*�ʟ�0u�1��48����م=N��|��.����P@��	����
������FzWӸ���b��J�]��N�z�In�S!��Ե\��͞YS�=����n��u�p��Rm��lX*�(����a���؋�~]�yT`�/�1�TK����������=�� �K>c3�(�������+�W� n�ϑ!��48zF�����2�l�fh����c-�S�k��*
"=����/�xˈ���4�`�\ٺ�E�x߇+���٪��O�ӟJwX����9�Ң�(?��m��d�W)�t���/�+�,l��f�͘0SR�ER�eb ��6�ς/�~����X}o{��?�C����9�.8���n�Қ��5�ư�jg�s`�"���TV��C��$gh|R�"�G精��J�����CD(4�U�E�Z�o�_h��0y��jo��r�;�����^�/�5�z�MLқ�wh�}���z�Gk���6�;��Z��k��7\��$�n7�Yp������y:f(S���S��_z���}mBXCՒ�Wlt���ڠH$�CO��G� ���Bz�#����_Y�#������x@?uњ���M�;ʚ(��n4ĕOv$@��@u�MZ��Uh��{� \����򱚕	ӷ/�V�� ��PXn���|��1�I���U�t�\O!��\EG�`�lD
�aV�ѡJ��rE'�V��&�2G�J	Ȗ�jq�[������N���>�W�X�� ?�I�*�e�M���N���d�F�^���?�Q�H���l	q��Q��(y!E�cu	О���h�����K媂�ҧ�2e ��D\���D�����I��Dp���Jyz�>;["'+O�v\J=늰��26j��}vM������3�vBfWA�2���F⼨(��xvmd?��3�:�u�9�LG-=����\O`4S}eiK��a�Wz��u�:Z>�ILnփ����a�	4d�U��> �n'�%�8͟u��lp^ �]���a�d�6������' �<��^�HC���`�"xP�����7Z>�\s��їb��M ��E�f�B�硌}Nq:�^�`#3��������e�{���7 ?:�؋ʧR�JY��h��`Bbg�-��2���c���Zʔݣj(ɒ��;}B͆��"��`�!���o�A/E��r6LܔX����1oW���y4�����&{;N�"���̕��t�IL9��[j N2��S��OL�~v4�̓����k�M;N,@�U�ʦXC��Ę8���+�_0�N����~(X~bXW�M*"��bbZ5�����(ː�O�	��0Q�v���#ssy����xĬSJ8�h�K��G��AT$�K���=�z�U�T���=�w �	9���-�����1����]��wH�	)�My��D%��x�9����s)L�,��{��n!�f^���y�= ��@�2�暎����{�Eo���q�JS;��u `�G�����Ә�r�[��+��@T]�;~�'I0�%jHf�X�#��EiNL�?�g�4���FRu�Y�h�s��M�_���ܵ����n79u�����֡��4�7� ������g.�b��E�Q2� >��K��~�]���5�����k��BOwg��S=~�6� n��i���9��W���?t���0*i�K�z��^/�M�%������7-�]B՘�u�e�J�VE��#���'�<.+�ox�5yo��l�����Ed_��h)hÌ����]�)ƱJ1	h����2�
D��ݝ%�.��z�B��.'����.d��?ϕ�K��*���G�Z���l���qL�Eܾu������|M���ȝ�8��KX��/����l�T��6���Zh�0!B��'�i{��I�!$T�5����&�O�6�cj���>ȗ��G�u�t�2/�5�m�4�(B���L{t�2�5/�ʏ��F����V�4��vtC���*�]}��Y�s�ǈ��|V�@�;������Nb��So������v/;�b��ƶ.�U�-��_Y�����!:���c�������v�\���x�''�*�����	q±hŮm��n�&y��!��f]�վ�l�X&Y�'k�ǭ����#?YT��A���}�8�=��Ys��Qo��Kw��x���&f�]�H���;��u�߳N�lLr���n'�L�&������|^�bʕ]����cy%61���q����_�$������B���D9�G��3k?�P��cg��8�-��:�\�m�Ȕ+���̉ �5�^�ɱ��䃼aգ+��֊�2d�C����[|�ѷV�Ԡ��!&��@o���;[DD.�b{.ƽ�.Z���v�~9+Y���*���6��a�S~�#�+3��$/�}�7lu�Q�n񹘌>3�GxWc�T�c��<���Dݓ�~Љ´�n���3�U_ɺK��iT���wi#��y�P�m��]�%W��|�gj�� t^�ߋ�2ݧ����=�V+R؁
�
|�,�eʵVi+���wd�V�p�G��mD�l>��1"�]����Ax����҆Eax�%�N��F���[����NO@��O�wq~�L&G��y���*��efBd����S9Dp��燻L�o��(G��킅8{,�f�s$�B�k'v3&6./z9�H@7
� �|�,�d��4	?�3#�`�)vHl0i�Z=���][)�-M���H+P.�JS�J�H_��ʏ��ȷ;3MM#���5�/X�ܠt�#k�ale�H�p~sTʖ9���n�Js�H���Ux�^���win*_����g*|ۄ�`"�S�9Γ�Q��N���\_�������7���4Qf4�dA�n�cjjq��StA� �Gr��{σM@�4Ӡ�褧b�����|	[���A��|�'�)�YĲ�����`����I��ٖ����_��ȋ��?�$�Y�N)�A~&��&��w3͏0�Rd��)�	9��دlk��I.���ٽgM	�M�����n�U�Q���U.?C�n{θ`�r�߃���P�P��8'���תּCt��q~���M½��Y����|K�:��@ȿ�hv���p��_>�Gnw�@Բ5���PwRH�n��nn�����v.�i\��Xa��a�x��f�1�z6ALX�~|�Ťk����.U��b����E��|�t�5�����آ�?�q'�$�W��]w 45��(4�o��,�@E���UL<���a�Wf��ld�QF}UF�c����G���W���ȣ`���:�G;��[�nh��U��R���J��j�i	Cp������:~�`�^X7ꓵz���r[�X�v����������[l#�p�)I����]���-���_�r�BH�=x����w�Xz��S1�l|7�kEs/}������
Ѵ���' N���3;�%U�Y*��S��j0 He�O��V�r�(�&y&y{!d��<�淞��W;(�d�U����uбOF�J54�*~I�B��!���T��3���?���LZ߅�l2����1ݵ�&��	-���`��l�M� �
�{"�/D���j��<��N�^�p�h���sk��8�p���nB)\U�H�F��ŨČ�=e��y�ւ!HX�4P+����"���<e��%6��$\�'������{�uǻ�f��wY�\�Y�V^24���z��j�X;DF�FHA�ybۑ?�I�%,��-���y�!�0�;`�����?A#XT�L�m���V����]u��[u�:���r���L=�DŊ�>�}�VZՃf����P4�gvue{1 Ll;��7�Ԙ%��#J��3�R۹S-�%�+��ө�ŀj<P�'Ku��H��lp�/�%F�o����y�;0{�Xu)��9>�pכd���_" �,��h:S�y|"�5azt�H0(��3�W0i��,)`��Ʉ�[�Ο���X>uR��8&�Ɵ�y�m3UGĘSQ���҅w�y�����K E�m�f����j�d>)�mb(���w�a�3��`��ا��mũ�+֩�*���9�d�5��Jg����x����<BSHp��n Mbt������d�L���-�
�g ~���Pҡ ��2�c�j92�>$��y�����Z�?������uWX�ϫJ�;��C�C��0�������+��G"j����$_�"1�C�� ���cN
�/��[��1��W.v}�5���;ۖJɥќ��T�dh�p�Ms]=H-� ��ؼ���Q W��};��\�*^Q�Ͷ��wߔRs#>n�S�t�!r����]�O,�E	SC�kE�D^��A�^��V1@��F�M�^󌏹�g����oeZQ�q�<`/ km�|���>�=��z�c��lI�P��گ#H���`�)xIn[oܷDdP_��ʑƮ��_3^8���H���N��W��V���˺�;8C�;VW��|�uՌ��>�t`�ӛ����HcV6�!������������5Y�Ƹ�rq�Ť��a\������٬3��{����ߨU��<���)�����l$gr��w��
?b�T��G��ZF�<��k���ky�8��`���x�
p(�*"�[[\ƫ�JN���b�4N���!�A1W�BN3��ҷ��bUI�Ub���ځ4�G�ެ�h�gZp$Ө+����_2��UplG�{������.Y����߼:�T6���j�鼜B�>��ԏ�!�ܩ.�H��_���|�����;�,_9��&��>HF�������ӈF� O�;7���aP"[乃�����En��+o��U�T	e��FE������1��tw����Ev\��o徤�y�����Q*S�	�R~Gd��U�xA/�"��g���Sc�ƕ=P�;+
0	����w��1�%�NL����ҼZ�瘝5o��s%CO١���� [�)��Ա�[��2�Ge�\�"���旿^!\n��d�|0����WO��4�.�@�lG���j�t�]�����(D</��`��g���Y*![��|	Hr`&<;�wB�M!�V�f��$������RL�M� ����Y��v�ewld����^�����\�A_�n����vv�NY6l�.X�/4�%T�9�奈�`:�jt�FiL�R�O�v��