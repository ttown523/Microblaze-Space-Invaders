XlxV64EB    88b3    1c00�D�k��w�Ro{Ş��� +^�A+x�����ؑU����q�T����|���m��eI�C���2�_O�.͜<7���zAnRy��AH@MDl|��\{8�!�~���	�=�δ]y���$e��� �O�X&�1:���� ��w�Jn�6���*4�C:�`�ڽ#��_�d�����3x{t�9��c�{oq�m�1Y�D�8���0��h�͕�j�ħ�Ɲ��d�J
��ԽMBg�yHn>%Ɨ�j�Q���/gK�C���~ʊ�	��� ^�ut�<��aH�y	�����p�1_�8��8|=� .-�v�]���1#$��"�,X2�I�r��-��1J��s/�^�} I�A�xh��U�>��[ �l���"M2�c�럑��hm�
՝T;m��0�[�;�vpCÞ�����r�e������C�*�X	CV{�K�blO `C����� ؙ��<χ��Z_?:Ew�H��5�j�c���o5���@��0����	�A�.к�ڪ������)��	�g�t�
�86
�e�Db��-~���b.��ͧ���܎��	��u�*�n]��%�	Ƶ���4����	���ƙYx��"a�����64V@��Tv��t�O������*��l��.��}�	$�W�I�m39�(�uPP��W.�<FE����W$�3)��7��|��xi�lLz�B{�+��KFʂ�B�l:G�v>*1���70�j�D?��HX�49�HG�����Z3�,��1;�i��&�\=���b/���&��%M���ڑ�4�6�'S�P�.�OAy���.�ɓ{
>j�H����͂+��/i��`�?P�C]��$�X�=Ͳ�YFTտS�z�l��TЊ)g��O�MG�@�i��,1�p�ŮRi��]J�7��ʪ �)��>�ȩ����|_D6��M��>L#�P4@�~(�o��b �t�:���ʀ���lBxe7���m2��+��b��ĵ�"A৏ )$����0�0�����%�u ��VN�UJ�>7� ��!Uڛ �1�w��]z�����ga\1��'W�QnJ��xO7��%)���ڃ�{�Q$�����	���2+�'�˙�aj+6.�L��ܝ`�-�k��xGHN?��7pAx�#o��A)���ص�w<�r���{�l�9�2&
񥗘3Z6=�y�f�~~��e��p�CA���L~Ӊf�f��������ȗJBC����l�)YL��l�:��B�,���V��s��3Ǵ���#��+K�b�q�oӥ�o��j�� �����-j�J��Σ���
�Vg�GWy��+ܚ�L"�z��m��8�w����S�u����v��#��+���v! �\���ߖ�\�F�'�G�t��|��IJ��wO�����OǬ�a��N�/D1���A����ˮ�5�XB�e��ο��������.��0����D�wυ�gg�(���=�pW(����L�
�f<���ie=��li����Xt~O����?ɪߑz��/ϳ >38Ӝ���=:<O=��\?[>87��牨N���Mn�C��-�h�'������-צk�+1&F��`V@��ug��+慬o��O�[�=��D��vd����+�|�������{ȋ����(�oK�9 B�4i���~q��,��ɓ�`c��,P��i'����n(�+��B����,�@�m5���}��񖩳:u�II�O�����d�����5�$��=K�/��%�v4���K�m\�]-��FF�����-�U(��1v��u<�@���Yz$�*�Cx,T���
�^�Z���L�l<��D\�3���G�!������F&�i���sVR޲y"�DFWô)W��1�zV[�����G���+(^�͵�	�}s6$;p��V�V����5D��Ü5��*��:��H�V�!q�?�E{[�U�Jk�Ϯ4��"�Z�ґP���%���W"��xº�\�>C�8�w@� �ӫ����h��f�ǡ�W�sp�|�:���̝�G�!�����o�[�H>#��l��A�����ɹCe �yN�7���n�R���Y8L�x���jJ��-�b��骒��o��`�1����RD)��47C�3��М�A��z�z�UZmr�_�-�,����%Y�QiM �{P��2��D5���c(R8oFG�	����^!3n���:�I����֑$�����!X�	�d�n�[<{�1#Jq�=Z�*�m�G0�֖A���6���[����%����4��D�����@�j�6�rD9LP�
"�a�ڀ&����*h�~�U�J��:e����?ɜIMXWB�8�Sy�C��*�.�����Dd\�YBS'�d,Xb��o���Wf��@9��:�N��V��N�ޑ�o⤓�y׀�Q�t�P�ө� ��#��V��۹���c�C�ʰ��s���*�W�w���މ4��#-�~B�?��!u���-��"�>�z�oq���!����L�V뚘��q��i���j�OQ��J���2m �«W�d�qv�Ti5�:0��(9��,�f� 0N�X�f�k{����p��|O�d�@t���C�b&h���?�^�}�9�;�p���ky���u�N��y`��U������P��t�a��Us� ��c|%�� �tp�&��uZ=O=��I�5�(��zc��1Am'�g8��l���tl����
�pW�\2�c�(���,]����� Y�A~��fi7]�e<H�{ �A���eBa�	'�Ƙ��|�|��&�n���ך����o��
VU��+De�V��Ȑ5׷×�YQ�y�/������O�����\ �K����I��6��K:�Ҥ�՞����hv+a����<�����Tܽ7%l��S:�?���}u�n&�"����)sHu�\�Ǐ`�Jv�u6�Ry�P{�Bs��[fۤ_ք�K�Ϝ���PuM3���!������R��Z?���(V:C�@m�3�����Nq$~�y,�R��7]�]"���Gz}���\w�� ��&��Ν~��7�s���6P�K��z��K���6r
�iN�B��X!�q8�}5^���Iz�p�G�vG��#E0�I�m�� y�8� �QM#�i��ݖI�s�,���]<L�����T�.�]=�G�WY0DJg���oi>3���U�<���L9N��-�f@�t7����ҧ<	m�v�,��U�ˏN�~x���%��x'�y���<�Y1鵛\f�c�/�n��!f�vȴ�F��h=8�p�y�0������;xJ�E	>F)�ب�#��Q(���T��[C&
�?��T��듭L�^���'���~s�ٷ��=W_�`/���.�Yf�K��ֹݨV[��~�#��@�'�H�w4g"��*NN����р�t�8ދ�by!�4�b�dg��Y�pI�ꜮB�'*b��*%�
��������j*V�OM\����ӓj/.�4ؠ-�:2V��RROȽ��)N��~�;�zm�fD�������X�$,���8�g���'H[�wp�>A��?�t6��BW �ha#+�iGQ����������ɵˌ!�*�)����>;o�SЯq9Io�Տ�x�?�n��g\Y0Qr������ ��O3���&c�sa�$�L^T�:�M�:' �'H/�+Bm �¨d���D�=�&�č7��o��X:��]�{����|��qh��er#���?�&lp��j�9���"g�)�r����H��֣α+y]�Aнuh�@���p|~_�B7�k�M+���Cs�`�2���S�>��<�Å�F�a�Pݦ ��Xĥ¶��;�L�^�6,f�g'�p��;�ͽ5��eb�2��[/
�3a��ƺ��3��Th�� �s��=���MmDS2#QOX��O�{*#�#�����fCى�2lz41L��ެ11C�|Jk��9=*���"�/0Gp�E��@U�6/��/P�V��:#٫���"7�9��p>���1D���,M��U݇q���'б䎀�̦�mez�u�Ty��q�Šh�R��5��Q�@�*S&��ׇI[�g�	��s��_�ǁ�V�*D��Y"�mNe3���l^FjO_�,8G�.,*p���� b�,�O�O`~�oI@���,gֿB$�����C�d$��'�?n�YU�2�-:E�_�׃	�[���rg�	p�+RL <�0.�����_f��<�4��ƿQ+nS"�eO��W�^3zM3Su�DK���Lsb)t|�V�:#�׌U-#��X{��|�=G���VR�\g!�u6�Q*�<]E�} �e��Ó����w#�x���3��$��Q��B!S�I��`���殁������8X�Dű`k���;#-�n�A�2��j��G3����Y�k��i5g��WW��mɱ.>\��ː��B���옃�f-WQv�ѷe�l��m���3D��Z3��7K�?~�L�oj��C|��f����˥2x��k�z���mg@�\��<��i\��A�������l�� xs��݄�VT�u:1y�E���k��4]�3� W_ޮ���j|!�����C��RM�wz�&�=3��5b�T[UcWG��f���rsźRD;�>�ݤ.��_��6�dlp�wZ5��T����͔�t���.K��bEF�]��ĈC�\㇌Z�ٗ�ɨ}*��s�hwE��ww�"��$y̐]��*�՛X��#�jU���IA�;�ь`�o�T�8xl�ko��&%�Y~�D,�ɱ��Ӷɪ:�r8�y��\����d�ӻ�9K�yy�˽p�A%R��DJ�����_L{}d�X�[��n2d��n�F��d�E�Q_����?�w����0����NE��dr@[
�^��~f��ÿ�U�hD�Q
Y�`�A6v�g��+OF��1�=.���F��Ͳ)�-F-�W�����%j�|r.�r�2[�6�����/O���0��+��Ў�6�Ĝxc��.6�ԁ�ܳt��3Ff@}S�[Xf��3	p��j�K ���F}m�W������+mj|֩#����}X�vҜQ�޽��(��c�p�Zoң�.G�������}�QKܫM�g!p3�&C�y<ćɸH��}���Kk!>���I]�����qQJ���3�?����/�"�I�u.�O�jJCs�HbH0bM��j%�u���z��W�ۖ ��ζΤά�M�k��b����`��FD��vJ����JE�1�$r^%Ӹ��	|�������,����"�LT1�m�SP������}�^�,p�5D�Q�u[��V~V�,�����HƢd(t����W�A�T_^7���H*��K�/��z/�Wvfg�H\�i*��"W�H�|O���$5�@�ʩH&�_��@2a��?�B^�~�m|ь g�}����Ea\��V��<�->���DS��h�-�Oo	uu^T!�6�V�Y;_d2j@/.�8cu��W�XV�ٌO8�*���\�v�!����:.V�ai��絛�ni^z+���-�>���>E6F5�Lo".1�6��������tT�;w=�X�
��,�J-Ʊ�f�p�����%�3o��٘�8ZâqT����eӛ% ��;>�%�N(�L�>�?���dD�<b	�eɛ�ރ�C旝]ZdID�҆�^X_	��f5R��oE����j\�6ZƯ��H�Ҫ;���(���ͺ`�K]X�vz��}�	��r���\�A�O�@7���"��LR�a3	�1��O���H���ܿ(�5ų4��ҨHex't��dp����4�_���~�W�e/���uN��=���0��&~z��Q���IZ���}��C^}F��������G1��X1����V�я�߯�
�'_��G._\i�/��%3/�et��DDd�����.�Єz	���>����:�w��)߅qU�p%��nJ��^x`�鮲~��P�T�k�!Q��93���k$u>󦳳��/O~��b��jm�	X-g�������3E�чw��k�d�`|���F�;,1�<����q�3���]��,ְ�c%���n���;x%�+A�i��}�g���i�D��D;��UR!��P�U�#Fi���7 ���s��o�G�e�0������qBV����T��ڰ�lO�먌�ۄ��B�J���Ò�Lޟs���70ӞS�$LFy�X�;��u<*߆(Y����E|[�?10g���x�f�����x������PuYHx�:B;�q�2�F�¾�B���!������yY���}�C�6�E*z�j���$�i��H�F��m���g��Ŵa�&��`����	d�]�W���(+./�g��T~�ҟI$��G����'�`o�*48���3�22�!H�u�\Y���kc�:�J��Q��#��M�X0�~]�܀S�����2�F���yw��/e��	d�ks��8�*��9
'��J�T��~&�u�1�[�y�]U���ZxK��۵�"˕����F���!ɿq��ݦ�S�u��T���J��	NCwe�ḭ��k˳j���_����c�Q/�<N̹�^рakT.-|�lH*�0��<���] ��m�kPi�>�o��r��nxsNg8�O��v�J�"ݑ#�����^V�}�[��	^/�ɔ/�T4w�"̓�E��W32���PE��@�m$L����H���₂]�eE�f{]&��$�L�>��V��i�#�?�l=�>D<��ェ�µ�7�v^�\<xQ��L
>�"J�j~��)�̞_���;,���|�Xn��9�B.��rP@���;%��W�kh��&m�$�S
2\o���v�y�FF�G$�����%r;���Ҭ�,O$�+ NS1�5;d�K��'	�qiL	$a^�K��f�\�?��X��Mb8H@h�=���E2}X�U�n�"S�Ӧ;�e����(����+����\ݹu�y�f>b�&�WxP�