XlxV64EB    56da    1340�"]z:)iv��B�YQ[��zRV���=qk�c0jÆs�D��������fJŲ(Oja��k�0��t�F��5��5����6����ĉeJ*J8�G��s���M�H�A�,�����#�+Zb��@�v��]`���+��\6[cd;����[�;���iw4�B�������*_I=1{�U2�����a��<{L:k)�s,��l|PL.�Q�e��Y���a����*�����O�|~���a�F5�w�r5������њ���#���݆�6=�P�xpp
�W�@����������)����o��OAx��O��,G�3��+�^�x8�%6����,XJs`��o�v똀�{y�<���,�&i�r-�G�Й��I,�PcI vg8�(���TgP����K�j�h�!<��ǡ��ҧ�Y�'<���Y����O���3�k"M*~�%��&C�&>����%J8��J��ܕ7�zb����-"�	2l�������\�2$'�5-lX�,`�����H�eB2�ߢ<>�E�
HAa'/�x�I��c@��z8��RÚ0�3�.@0���^bKK�.�6.�c�S������5P/�5yQs�3ó���&T@򫧼9�R�k)�qe�X�S��"����9>��b�>?��T�5{r��W:�r-��Ŕ�򤲇n$�B�|xo�b5}�T��-??S�̫��o>jrl�H�. ��ʟ�C'�5���j�o]?.���v��H�g&�.)�/�l����>H+����8z[~"���x��=����:V"�K��(����z�OfG�F�gJ���R�H�4V(C>�/��6�6,ɠ���eI@!�C�f��{��2�M]��%b;��52�y���7��Y�t��F,ܦ"��ǅn�YP�o���1J���L�wZHt�>]�o��;1ٌW�W����:��a��L���gj��~$ʋ��{W< b�@��7��*�/Ik�h*]l�"�R�:��0�(|jPɡ��g��닾fbt�y��Ol{�8�)��c��33D��0~����_h��$�;+��yp��$����j����c� T�������'�֎n�o^���{[�`D��0�~�nOM	�t��|w�7�.�)n|�3�)����!�A�$[�kJR
j��3�c:�d��t��ˆʐTM�T�]�h�/:��[�J���|+��l��7�j`Ms���5�ә��:�%7�x-K�kT6�����)�;^w@���5�<V�ء��,�PU��+~�w�]��)i���Q�ވx�OU櫕Z�b�S��Kp�G�Q��ڮ���?�W3�)8�S���~�N��ܫ��/4�[E���v�P����`a;k��o«��6��9�eN��׶9�[;��F��T��_���PO.M*E�< ���U��Ɋe����[�h��tʳ����_7��tnҊ�
�,���-��n:�c�qͱ� �s0�ۧ~$ ꭟ;43�r����
�����NT��i���u� x��ă=|��v�&��7VZw�݈}�˛	�g-i=�
��m�S�u�6q/�z�����,�m�\0ðxe3��.-s�b)G�����oE)�B.�M�|":,<Z��y��h�*�xx1��B�u�����kz��l�Ἕ��th9��)��1f��ܳt��wL�PU�7t<�h	�QN�V�J�������@��UBP�gP�4���>��U�j+٢�)H��Kل��F���Ո��Ɉ<w�ɖ2�|x�n ���5H�˯�t��s���Z�j�c������#�:7[,&��'��}��I����lh���mAk�[	C�ve�O1����9�>�{A"Ƕ�2�aZ@��RÍF��[�+̟X���վ]�sqӲ��/ޠ��
r�`� }��ْ�����L`aօ��<�xeJ~�U�wO5_�Σ���@���}�i<�2�ŶW��"�B*f����9ȼ���yd4g���j.,p?�%RZ�	�s���S�f�v�q4Ήv�������N�GL)T�3
���z�%��wpU戀�Kl�OE�zs
�J��)��|��\L�wAZ3i4:�c�� M\����_W�����wdgc�h�����el�P�g4�}]&*�ʜ{o:�������4v�?{aߠ)|-X7p�$ćf���8�P�즗":��g/�לc��m)��.ֲ}���0u�S"R��	IR.J�Kmn%���	VF�M�@[�b����4�D���S��$$"�
'���[A-�����S�����S_m+j�;�SH�i�.%�X��Q"��@� S�E1{p&���h�Z��%a�>���ݱ�6u.u�*'�u�5�2H8���ݯ���>�����n#����Y�`/�>�G.Gxw)�$���tw볞��lfz:����#�t�&�u�U�n�~,IA0t����	ezpf�N��d�܃?�S�I��6 ���?]���w옷�����d���Ѳ�pW����=݂^}`���.�ۖ��U���S�n0[�,�Y��V�%JV�WU��1~�V!��ƥi�|�C2� 6�1���ϬQ��^DI��b�n�?ʒm�gz�_"�����n�L	�k,+_
�y��B��V��t�\�U�g�z�MD�Ɏ]=8�R�'��@�T���R��NU_��hF=	��Ɲ�$G��N��<��6,2���Ih1��*��Ώ7rk׉���3��F4��a�FF�@�:�wz(-�n���x�4 �s*B������ᘋk�"�9X��B ,M~�Ʃ�C	�>Xv��m;�-�]ZW
f���A��R�㡶�B�`�3�����LU�<�I���c�e}LڳV֪5��S:̿[�x�V%?w��_J:e�SIH.�i�������UqP@�ڏ[��z��e����qV�%Ju|R݋�L�O���5���np�������@R��)@�[�㾲�PU?u^{�I�U�<�䲥�귰�M��z���j�
�j�`��,ۆk�PO}�9�cH�t���\7`>�Bf9�')	�o\�B�K�������m.���r'0^*Dv[�),��a�E�Z�2���^	�����o*�!a�DE�٨�%{/�XoY�*�G��U��V��
���G��<�gj�UJ9S�|^���wx����W�a���_?ńJM/�����[���Ե#�4�����/�)�+��V���j!�?����֠�Z�0a���TPh���&��I��Kq��o����d��Tʆ�o�_rx��X�\G����v���Û�F#u���t/�П��0�u�B`��0\��ݗ�p N�fj����n�9���k*I^�5����/q\Y����G��%��"�v�<iz���2)�vQȬ.b�őn�ۿ�^��j9�)U�B�"r���0��I��JU��ˋ&8k���
TEug����EE�'�W��U��o�Gm��hOfꜜa�7�2M=o��ɇ �Z=�)��t��}�s��\��FHχP��R�����UV/SE��b���hbSq+Q	Տ�g��	C���Jn��ĝ<�e���{.�WI?WL�Uqp"�͐5���n~�F��M[��q��نm�hL.Q���x��Y�P�!��< ��$��M}ȟ�u��z	���Řy �A;Κ����h��{Ƣ#�'oޑ�z�&��E��Wi5�F1��#����ON����e!l'�Q����9����J�I� B�aiy�AueD�0�0����6ςs�2�ݕ��ɨ�/"a�p
)�'���H�ƙH]b���f��O�d��xN�_�j}E9����
�UP�9w�~�>�<#̵[�?�y��i@v2g�P�sg>W@�ՙu���RQ��T�+�ա�
a�	�i��A�1��Վ/�Z����?3M��u
�ȫ��gT�@�7v�'� �+f�5���H�8���LztB��GH�����߃���qF�т�z�C��$��S��xZ�5�5�	��F�K	P)�=w�P$�>R�鈇�2 �i���:��+n)�8��]k��smQ�������V�� h�t�i�͡�/v���J�'?���|���{4�Q�N9�iى9Z��u�G8x����}I͆������CضȮi�i�Du6�'�Zu�%鑯�[6q��Rd�����'R�����Ty��|S>C�)�[~v��C�H}�F�<<�tfu�?>�&�;��g� �繰�/���?���c�,Ȩ}� 9��\��ۺx��W����o�m�����C� ��C��1O�D�T&��h⭑DNb~d3�y�g���.$f���Q_,��n�	��-��\�LbA�չ:�w�h�1�V��\��ޞ����|" � ��u�0O)2������n=�q��JPtAoS�0�C�7+�h<��2��/��y�%�T���U�x�-F�Z�!�1�a I �ր��buc������=���q�����D���٦|t����{0'�v$p(�A��+�o��O�3����$��N�1v����y�!�A����4D.�%Ȼ�ςI۴	�(*�	��?��5ǘU���Z���lS�T�h���_�R�0M[	���ʙ�
�W6���u/ ��<q�zgb���,�ݕ�J��]�mt��@�����?��z��#�$��'��\Z�ĥSc�kW@�(�nG�5pΞ\'�Hf��~oi�6=�"NX���	Z�Icd�^�m����� ��Vd��on�~��"��hW^Y�Ǳ��,��/;��������U��1�{�=�w{2��]ɥ)�w�p	�D%��^�!���K�E��	ܒ�M�u�=�*��