XlxV64EB    fa00    2310���ħ�f3?p�2L6e'�t�c.)���N���9���"��u���a=���S�ه���� 7_%1�����؄�%汧"����>i���#�"��$��O�܏h����"��H����C��5�(S\�DA0�c��&�i�K�d2 �KO���PO�h��ffi� 5��T�`��a�&�]A������j$��S3��_�B���,"	!v&4��{:�Y>��wD��"{�ӷq�mC���q?���i�B��0�yJ`:�0Z�yR4�Sy{��P
�,l�b��^o����$$��2Ѯl�3�NI�������7�K_)���B!2̹A ��D���i�%Ҋ�6fB�����CO��t����_������ٿi�����R�&�����)�M�}Nu�VĮ.��~chd�����o��T�,�@��B�ΪS�5h��u���#_���IO���� ���'���a��9�������ۈ�"�׀��<�ɮ�W���a���[�̷���F�aJ��w�v�����$�YG���|��˼C�������
c�����Z�Y߅��+j�
t;-���pw%gw�d,'���R�L�����촧 �`�'����Il�Ϭ]E_�/#3ķ�q�
�ڳ���qR�B�w�S~�g
p�RE�12�)j�is"z��E	��� ������S�io�7��Jv���,{��#����p�;�;��7��M�p4���z	��5*�B̖߲ݑ��w�B����5P�ߤ��&v���DV��W�~ST��b�􂟫��hR�LȒ�M\b'��.��0�B�h���;toU��.�1�XB��"��`�i��L<�O���r�,Z��[�*J��1V>��+aRgiZ?:=Hj�8j04R �.����䒩�*�BuѪܾc�A��|ގ֚9��P�u�v�X��[��ʠ�\�9"0>�^}��|sSJ���uo���:�b65`��%OF�w�؍&�]��a��8?��J!��Ҋ��=�$��a�r����lU�j~��l�C����.���T���"����O�2ʷ��<p?��x�d�u�~$DX5A#oc����2�A�@}a�j�*�h��B��?ެ̶�~��8��ė���a���oh�UT��!�;T��]v��-Zv�\x��N���Q�p�ʉ�NN�r)���~n����s^q�G�NT����o���o������ٶ�q"�hc���7� (~7G)ʃ4l���#P������Rc�?�~K���6�P-y��ѱ��
�eN°UM����� GWg�D�f��qS�<�HHT�I����f���Ӄ=�� ����e�4�FF �-EȚ\X��$��=b��9��@����̝�^D����`�x�����T����$��"Lc�]mȀb���.Ӷ�l"�}uT&B�k4VIye�OƏ�pጧ�G���ذ�U�w"ፗ���W��N��FD|��wf_��t���u�Q��n�P�)�:� �!���ٝ��s�z�5.y����"��l�olϡ!i�_+�J0�p4� ��Z��
���'#6�`��CvڬTH�����I@����~�`��fl�Hg�~�_�R1e��#�Q��L~����A�n3�"�(4dL�������T���0�,����Z�P0e&�i��P�u�WLh^~�j\�$O���0|
�T��*�Sĉ�����C�H� �A��e�������H���}���Y�V�O⪣��b�~v1y�s��]O��k}��G��3�͛*�1`�w��n-�dz�=��0껀P2�[Ȧ����
�+
h
Boyq����s7�tx�!��_�_]CK9���R�:�sfh���guO#�>=v��� ��G^��Qj�c�����9�K�a\��U�Y��T�~��/F��'Z.�%y~B�_�X��R,��gP�2���� ��«b�pԡʇ�����dH���VT���}x���G[���S��t_��ݯF�i���&���a��΂�7���D�������V}�%����́���ZRn��c�Ԡ�����-d�5����%���u`�{�Hu¨��@�Y#�a�xX���d����.&�t�����	�o!è(­}Sx�D7�p���E\��ҿ?�u<������G�+�6�^oa^�Ӊ���6
�0�o�����+Y�U�^�+I�$���xh��e�V"�����04��_��o��c��Cp\�GD5Ruo��ט��j��@m>��>XT��!	�:����\�	��
�c��6�U�5Ŋ���nLf�9��Q���	��uR�������{x'Ys�=��%�8UJ+~�I[���"<֪�l���P��$ �S�{}�4�xEwA$��W�#��$��َ(%��u��^DuJ-�W�H��<�e[��s<��R������ӄ�4��g%�~�����`���|�?�ԟ�/弍������ �.P$vt�VG�2�b��/�$���NP<��h��s5���^H��c�O�/10����>��S�NX�ځ��Jkk�hY��-���<h!~�Af>	`�xe�̟���5�J�N�4��]N�Lt�O���lFE�	�1�i3���ߊaD���A߄���ۿ>�Cz�*�����@/|ޡ!:c+�C)�[`�`2C�j�4�����.��1)���V^�jx�_����3c�p	[apo�>ɽ�a���sA�? ��9(�^[��0�w�:�7��a�����0���ZEȇ�d��e��A�:u��N����[�F؄pf��eA\��Y%h�P`K2�����=�|]���gOb�>����UN��@���_]�Q�]>\��j�z�6G�MRH�b���;�%s$��ɡx��\�.�P(��<M���W�C����������b��(+Ē�&�!��n�Wgï�"��*����)��qc�r�2"�$��d��t���j�9-�?
�AQ��k�;���쎹C8rE�K�����e��3X��Mm�o1-�U��d[�4�%K��M������5�FRS��#�c�$�sԺ?��V�-�q��I����idޠx���p��ǌ�{)I}���ʚٕp��)�N�EaF�L�F��J�E�$��� =�$hQ���A�$͜���:�V?�zp>R�]�\�-�U�
P���o1
�
UX�y�p�h��um�yT�JO����(��"K�kb��74q��j�D8;��8���d� P����ۈ#�Ǯ3���Ɓ���:͍'������N�cy��Ɯ��Eb�=.�D��v(]Q�u��3#Ț��͏G�tM��Ӊ���{���M�T�����D������a֛�Y����lX���S\�t�m���Lߋ͜�@O�<h�٧166+vr�=Е��S��.v��:[i�n��W�Q��nX���M���fC�Jr&�W��"cfs��	_���
�h���n��tL��B�q�΂�su%_�����<�D�\�l�)ҟ�L����J�Gm	��%gHU����A9�c�1ZnpqcKօ�)Q��Z�O���DA/��	�� O���)�Uȯ�K��t���_P�7�fʳ_�~w�
���@��oDk.�-Ze�@7���O�;�%���q���s��D�F�<����̩�%��}
�t��`��?���p&�{p��%���r�ƨ�tx�MSפ�[���Փ�M�1�,��KӚqk�I�0s�kp�!ҔSROR���j��{?�`<���:!:gY�|��0�RV��W�	vٖ�`O�B��M)^�'J� ��K��ǭ�ؐ�Wr���!�7����vm7��h��(fi�_���w��},�k{�
��:k�LG���y,�f�~�Ik��7�\B=C�1�U�p3�
t��;��p�]ر����J���)���(˧��h|M�Z�t��;">Ie�ܖ>_����d2R���PZ�7��� ��\����^��耑�L������&��)�����H����$b�ïT��fI���'|z�e�3��+�i�J���)�t���yN�	x�ѯ2^��MC�����!w���@�6B#����`{z� KԫcNݦ�*���Dw���u�H�C��W�^C�I�z�'�j~tAջ}�+�cc�"6>7���6�ݛ+�&.i6%Ւ���J-��i4t	|OMYtXb��_Ӻ�2++���L0���_R�1�+6җl]+F�e�ꕳ�OG������wFӈe��BFZ�.d��g�#'��t&�o��a��lK�7�3]�f��=�<��K���Y���?�����0�R��)�_hhm�w�;~h�����KN�U�D�a�p����1.C��T�gd֌S��ژԄ��k͆n��>�B�		�Aq��A�YD!�{ �7k� ����Ј����̬�-�B1xȑ��[D�j瑪9�V�w�X`^�D��i�p�z����)2���;[T�N�-���AKXY��{M�AUHc��6��̘��E�yqF�*-����2<��S��	!$�i�w���\�[v��u�9tJk<���~1Ws<Egd�uV$�|G�Md�?E/�0f�ʹL�cE�g���K�s��`�2�~�Q	�����N�[{tPB�.]�.B�@3�l���Li�@��fX���ˀJ�t���_�n	(�.�^��}���:�}�HҖ��I�������P9��֐6(�>��-����	m�!m��|`������� wr�z|�}>4˝b�3������e��B���á����`���V��W�oI���:����E��' X��Aޑ��8(��zMҸ���o:��r�l �X˶F-8)p�<����ؿ�;�9,���*���h��L��Tk���X���#�L��[���W��!�9����3Q42q�@�p}��w��ٿ�����я|�c��Q��u����Y��V{�W ��/G����-|E�c��󚱌/5�c�I��F�t�(tu�Z)��qom��,5�v����_�ɚ#m�^��d�pc��IQ�BC�q�xEPaݱ����y>��(�Aqܝ��� �ӝ2S�A�`�F\:���K��,T����<�3ӈڅ���5���':��@FP�P�?v2Do��8��ر��,��mx�j�d¸?P�'��W��k�.�;T��k�a�=��(\|�?m�s�2�O#C;a�b�w�,�I)�a��h����-���P>n٫��Wf3^��]�O�HǜJu�+*�.?���.��}I�1�ݬ��B�������i���F�#�1Lߍr�ɦ��_���ΎDy5*�@�m�H�p�E	��t��WNo��Xw7L;�6Qb���U���w�uxwcu�CY�����)J~�x��8���k}s���l�"D�J �*��<^�p���
�p��\�^2�I0(���:����@��Ps%�Jhd���E���e��Ј#��Y߄e�J�{�^��/(����C� ��(L_H�e+�5CW�Z$d�uA��N2�wu�_@������J>2�Xh�|�оInw=�]�����Ǜ��$h �8��a\G�����B#}���//;��7�,�L%MT��ѻ��,\^���*��D��MM��o>Ryٓ��S{�M�K�_?0��f�]'}~IE=aCX�̐~cnO��͎�{�g#��euV�^��dU�o��؛�M��v������;�K�'��덏���1[?�m(6P�7��3g��8{��2����BmE��(!P�6}�k,���t>d��Ie���f4���9��*�i�����Q�QIO�͘x�4��,'�+�Y��@��Fބ��+7�7���a��L8ٵ�MN� ����eC�Mk�7n�����u=��-����BZ��j�5���	�}�t��J,/��9��Y��d+i!��F����e���gYA	݆k��������E������t&��Z���کw��vI�FJ����G�k�'Z �*�c��l��ă�0�S�e^��^�i�OXfI�>�{;$HJ�{�b,X�rg�ָP��R�h�#��B?������Y���L�-3!U�2x��/�{���b�l�Z�&�!L5Kv��� �;qsW	��Ҵ�w��z%�B?��m�s���JC�D�'��G�@�@���_���#���k��K1���\�6IR�����*w���!���Ň(��/?JG�b3d|_ѣ�N������E��i,�HH`��ş��
�9��EHҶ5��,�+����7�vIR�,�K ��}��-�$8�-�	=���$��>|�؜@��4�e����[�>�i_��2��Q��?@��O�ޟMh�Adc"6��_�-�����&�|���tq6Q��q���	��[J�ׂ{��-��,@��Yqh����N0%�iI��S��L��ⴈ���K���D��!5v���+h�456��Kl��jZ݀������ڴ�+ [�ٵ5��Eҏo�]�`r���<��ff��!>�MLv�-[�;�-(mɑ�x3��r.�y��x��wN=�}�է�/CB�R�	��T��	 �|y�WޢT��$�lV9�XBP���[�q��l���E}0�]�=�[��w���O���(6�щ 6�1[b�5�<E~j�S������ؚ����o��4�z�"��7Z�����
n�I �O7KJ�$p&�<��mNt�^��C�������QA��2��8����4�s�V�	,��n:�t��B8��y�Zi�vdej��Kи\�p@��̗,v��[�1�J�&�es3�X��*�2`{\��9�l�7��[���]���G��	� O���--i��e�@�'��#\W�O�g/�ZLL7�,�t��R\IJ���<&-燁VӺ#��Ёi�D�S�ʉV��3[;wjw[�e�	M�
+�[�~�_+��M��e�qS�s��2�0�)7��X�����������ǳ��"2I�l�a�w��tz�uXa�m�C�y�t�[�u-�c	�)�_�MQ�ߢ^��{�$J]%[x�L�ZD���?s�r:��8԰�~p�\IK�{���Hߟ��?vf�x�ݓ����,ݏ&y�נ���c��<��MKL�)#��X����c�I������<����G��-:Y<YF\$�	��L�f��
�6�h�O7�S�\�g���)�,?�������U���%��%��(��?q��\K��m��j�Y�6�a�'���+l{�~� Bj(7��_ϾT">�L���%g��?y�d�m�Z[gOjz��C6S�AV���#�6�t(�%E��e�Fv�br��p�	/�I��zq�9��AA+�{O:h��ej+��ql�͞�5`��Q�74�����e�VL*�bk��g����ͪ�|�X�&��@��+�w�fqk$0�h	���2�Â��:�Q&��}���{�O����w��sϰ@��.������a�?���C�Ɛ�B)C��c<vR��P}�e��䐹�l�O�eɯ��Ky~���7Av��郚�qc�����j�v��2��B$Ϲ��/�P�����x`"��(^�{���h�ʀ�c7AQ!�T �o���w�Y�����A:<؈`�}ԅ\Q���p<� ,�,�|F����o��W��IJ�VoXY�29��M���h=h��,�'� �m����T�іN��ZM�N<m�a��M�f���Oh`J#{��Ň�-ϷP<�K���p�}Ǜ�"�>
\ ���=�\;��;T�t��&dݓ�EU��C���m����1� �H�����؎���;IM�)���dy'@�v D�r�Qhù���LN99��W/O��-zC���N�u@+��Z��C��Ju>H� ?��]`���� �9!��I^�r�29+!z)<{�l.;1Oo���VgC��6dM�L�`�.�*љ�C/X��v��?�2�p�$�"O1�����#:?J���D>�9�r��;F�緰N���])<�B�2�9.��+�) �Yg�ĔA-�s��.�ap6AjA7�`��l�����9���|�ReN��li�F��tA%�oz�]��-����|J��jܣ��	�k*�P�@1
	4��Ft��KZ�Z�O��#�e���C
�sahb���T��)
��V��56)�R�d*)˺br;4���2w���E�dY�8�ͷ�~��+�V�3a|�7�3���#J`����x�-��φYm��I=��ݲf5fϑg�s�JS��F-?�m:�}OUp�E2�]/����G�1�_ P���\d����50�禤�V�,TS)�%��=��(�v|Ak���׸� �2�pÇ�QH���o��N@ʄ�M����#��x�Mɧ��j���}0iO������W�������ՠ�߰8���
�ӯ�P*�fl�V{��*���&@�������o=8uFZ* O�f|dV
�,g��y�de��L��}|�Q���Z8h�Pq����Ƌ���ji���'i���!��;�,���mt���z�ߣM]�p\�.�Ħ��,ᴕ��N��f�� m_c6]^�C
3�e��d1ZمA�ǽ��@��Bb2�x��\t�(2�:$Bx��9t�����rz�b3�����5�=���#�W�wOT	i�Dq
:�_�-L���B�L|�xE5:<lQ�FO����9ը�;�P�RҮ�6̣*�{�����NU'�|&R~���YT��;f�?T�;4�C�¸�;M2�$�V��g3Ƞ�2���O6���4�XָԜ��[�)
�]�����7vFWab)�Zy��t��X��bT""���#i���
�%�}#XlxV64EB    fa00    1770R��Rh���=��I���A��`��!k���� Ga|�=�ۡ���DMDc3��}Kx�]'��ZE��PȻ��/��Ոn��\��� �t�hs�",��ϕa�W���R#���g���8S5*�R��%�p!��$6�l�4����c�USV9�![��P8yQo:�X�|�D��S+H̰�j�4��D�0U�!��e��U�� ǀ��rk�?E�MD�~�|klg�����Gd�"txO/�?yW�M���)�[�%�������<�C����נ'i [�/�k<��f��[�Q1���q&iH�XQ���DG��m�Uc-��yJl�WLjX!6��_���қ/�Ge{�A8�Q��i�d�O�f���D��@�x/���C�I%��q�!�{��X ���� d�i���P���B�E��2J�/���clK!�{9��1I�_��֗)o��}l6ٌm��F��A� �C~I�D�4@A��a/���&�������po&�x�e)x:����}���f�S%��>ԢhR�?t�C�n��:��n�=�33$�u�����Ȱ�MV�t1(�� �����\�:B�a�[�:�#�������U�y�EiS�͡/��^��{le��r��s� ��}��G�h��Id�eqO$(�>[Y���c��C���ĥQ��� ���p[��)l�0�Y�f��6v�!��K���i���V
��a��."���1���i2E�Bb�(DJP2Ut��$ɹ��Z�9�M�����گ�|��;oX�!{2Ct61�ge���������#��!<���)��b,k�}��[Hu�ZR.�*4D��jJ�����`�[���Ӽe��D��m�d��a����	e�ܺA�g䀔���z�і�#2�]���ֲ+(>L�?�?v+=o��L��]Y�oݤ�3�}��o�A20��#+��G�e��{���)]�V��~M�(��9�Y���=�U�� ���+$��ċ�{$�Ӑ�����1�67�^�����!۾��_�u�m-��ޝ�5�y�y��>�
v�_evc���,�t-�&�O=W0�Y���J���=��ﳓ�9��A^��1��Rn��y�Oy���HM����@�;W�y��3`���e�,��t�0�/#�}�,wǷ��2͟�
����N�Ж�$��|J0���-�@W;4"qn�7�;��OA�/�5�>��$��k�J���c��=��2��c��-�7>�� �ڗ(D3��$ޱ��G�?$���
y�b�O�7��!��Ǚn�[�.��#DdI%���K��Ð�k�(�/Y�X]u0�,J��G��D ��H{�N��A�@����n �8�(���G�]���J�����K<�X��U�r3H�#����;*쌨�H%�K ΍x%Wb'�6����.g"�� �C�rH�*�6Sxì1���߃x��so�؊�6�nM�=����0� h��b�Ǣ����&A�q'�cY7ts��S9�����q�K�d0�������NK���mg��H��d[[�VI�6U���A�N�� ʧ��y|оs
�j]��#�M�� �n�*j᭯�z���mvA��YU�.��v/"e���Є&@AqmG�"���	A��~۝��g 95��h�}��D#��m���0��g�Z��ȸ�m�}'�[�6�����9|��X����`\3��ל������`H�C��c�ո�c��|a���e���nY���M�YJ�,Y��E!a�L����w%K�5�&Q�ak�\�}�
CC �K�΢�*��+\G:�0PH��g���w���d��2z�����B���d�x��yu%�7Jk^w�1�3�@���b�}1�l�D�y������k�Eu�f�&�d��z{�v�ĳq��^����I�z?�dWp������q�D�aRi�FZ�WK��R��6ǿ� [�)~y��?���;��뀋�O3Ƃ����'�bѲټ�jVj�)hj$���Ia^/q�fS�χ�hqZm�>0�c���\ZQ�i�+E�I>i��Ǣ���e�P$�.��0�r(X`Oɹ�"�Q�L��Σ��oo(�:�-m��x{#���ċ�Ȯ(�>�R�b��鸰��1��;�֔����X��b=G�Έ%F(�N��5��<,ټҳ��?gEZrt"D�L���zD\6jTO�ۨ��.��A ʏ��YG�X�h>����U��r�Q��e]�X�6��o�i�_d��ɾ��g���������Dn����[���}k#�V�Ҝ�0�C�j����	+�AQ�E���a~��
3t���� �#��P�5�ߜ�O������[�&�C��j?��dg���ָsjJ�s*� d���e7wc�.	(ɐ;�q
sc�}/�!�j�@:<����{eEʓ��ɕ��+`E�P���yg0~�.`�/I"^�46������Xy��<������n�U�W��#K��~�&�@��Y��k�v<�X-��/�dlq��
8�� �;��(����H�W8o!���

���J\ҽ~���@,iU���m<��P�Մ#�����
�;�.\5�ۜ����.KO��n���ps�J}B ���u�Ne�b��o�+�E�x�M�kdiU�?���{�*N��9�W>�t�U�)�M�֟P��P��/b��i��]n1��O	����	`������6�B'�]91U=�}���3ֽ��8�����W�[E�2�Ρ;&WiʮH���?}Le��L���~H�Jᴬ@�H��(���r^k��L��dmשի��}$y����R4i��#�'�8�$��k@��\#���ַ�����{�XW��M�^j�H��܎;����}��G����3cr�Զ���~N:n���R�>�B�q��剙j�@_'j��,K�kTC8}�%~�z&!8����q]&��1tr�p��VJf:Y��ÄP�Y�׼��j|5w��؟c���j�F�9ĝ4�6���M�j�������'f� ��\fk�hC�%�ۊ4&��F�(�M�X�7"���M$�erB
p�]��0��FvO�9��j� �.6(-t�� �2����"�bm�ʢ
� ��.b���:ԭ���xE:�&^}���^�͌�S�8����
�x�:��3i+lL�it9��6��tL؁��o~Z�-��4�J��|\������o"󹀉zb��no3)rT2��~]��<}K-����k�k�h/�f��g~��i7O�qU���v0�7k��T=�ُ�wP4y�>� �o�����H�AϚ�0��ʿ�Ֆ�����-i(;/����J=��(�I�l~0P4�^����Ӄ�zO1�ç��HG���W�^�����Z ��&L*�.��vp��/`O�-h�,�]P�/ ��sVB �>�SXO0�!wb�����~(��R�M����UL�kR�1���[+fj|
�[� z&�8-#d�dv�[��̰q���z �����:�&��<���������yt�� ���|����VG%�"����/��%VV�*�=�_��J������(��P���P��"�U�A٨a��1՚�.��޼��f�35��o�r�ό,~r3K�pץ
��E��^(��\2:ãn�S\������.�3*��r�_�ϥS�>�n�O/	"�{>��e(�������^<���Vmw����|'��7������\�a��u]�<֫�����	`>f��C
oٮh�C���M׻��H�kM�N����YOh�!��vƅZV?ItH�4��k�`�܅��Ⱛ �g�=i��m��|��{P��;�(F�	Is�b�(�2s�T��z{�z�xK����q�Tލ3��ބbB�@�Wj�}�p��q�A�������R�;�*�1�B�y	6X̓�{�P�]�,�(&O�)n������k(�>��f�.��;�0�(r�rn :���u�%ZR��7C�;эJݸV��>�)aO��		��H+7]
9֚Y�n,(s5�7ł+U���.6P�R�;�7I� x�?_w����y��$��븲7�H'o�e��ا�Z���d��y��2dI%`���@>	[JK�%z�Ү`u�Z�[nE}�d�)��T��qTW	�N�����1��`��`9MO�/�^�j40z��Y�kmƉ-�i���>;�4Eܰn<�/���#��9�FC��.5#��г$";���\�s�~��N���~hw���ט>��T�MVA��x�J��r�cyƱv�]��v�Z��Ǐ�绔����D�����椁1�s<X�[����� '�P��P��e��TE>9�8�E���u{��6��)��o��s�E�mR����� V���d~E����ԅ\>}��T4��yW�&&��ND�'�Xz�nka�<��>��m�I�{���jG��i����?�|q�yJ�M��c���Wg�"��!���x��ux���u�%9Wi���gɂ�җ�t�R����T��"��pTax4{�A��S��Ө/l��iX�Q���h�=:7s��*���e~����h/�
���k�ˢ ��[���A�V%�V������s�<�.�A<�吉\9p'OӒ��tl��M�u:�`�x����vZ	:	N��U�Rt�LO.�Î"쏵|�q����bcs�r)F�Fg�wf����XH��}�����a,[Ss�A�
�)������+��'�#��Pc�X[}�����&�è5���8e�u(RO���ZϨ)�8t���aJ�j�(e����ֆĉC��1��1S�qwn��E"���U��IJ��S��?a��[X��õ�\� r��h�����x���-�B�{�R�,��Y+�e�>Π0 !B���Q?Kz (�ӧ�{��y�6ɤ�h�����j�ͼ%�D����
�ⅈy�[�� �V�nB���y��>n �#��\=��s�7�JS^'�Z�VV�p�|�EO�=��I��p�y
.Q��g�z�5�ZYb�TE�w��������٭�ʎ��L���Vhg[a��[͛��g���<����5V�:��ͦP�b��MnZP+e]O��m�(�>��R���[����Q}� 4���p)V�/�Sr{��'(4��c@�?kU�����k��������C<��B\A)���%�2z�����k��_�_�t�S�xj��鰧�}.�%n��^ �d�0�ED�)̖��؅��|�EM�8x��l��a�	�jaQ��}��6�=�o���
�j��ۤ�[�W=��7l������2�DO�!Bfp��d���D�U
�5��~*'�K�^���iS�魎	w'�2M��1�Pv�#�ʞ��Md2>���}��06^��>����@ҝ���d`����S"2J��L��)�6�a��%�nj3m�Qw�楟ܴ
�� �_ra-K*�Xp�C��F���U���41Ң	^�R�s~���yY&�pp��e�F������d*;6���-r�#�M���9&����E�;c��ʠ��^I��=QP.J��^���мu�ab$|�;LOG�ڋ��������/PJ�T��m�[�)R�)��R&��J�hz%B,`S����|Y��&«IV���f��u b!0J�5�Qp[x�IϽV9���g��q��oe�!�a�o�zw�y���BΉ�Ho������=���+\�So�+�̦�.��q</��Eˊ�_��x�
�[�"�D�̄%:��E7��/�#O���f�R�Ycs�}��^�~�[����em$jy01��R�m�B�P?]�w�o'���>�?$���%�R��j���[L�r��K�t����*�|�܀t��:^B	6��s��Y���>\%[�zь�HϮ{S��AIQ�*s�g�i���16CXlxV64EB    fa00    1fa0z�	Dp������/u�qF\-�:-���:��$J��\�,���Hrs'��A, '�����4�����w:ʶ�tu����x*C(��7�Q�D�F)*����/�p���E�����v��+�=X&��t��x�x fV�&�^�g~ߖ�$p#Lb���>u�ba���h��C��y>P��ݫ��_':r3 "8 d�t��6xƧ��&_z������0T�}�M/߃āˊ�zno������d�D�D^Q�SA�e�diDg���@��8	�Y1B�rTsh�dw����ӿk���<���!��C�Q���u��G}�E��DX5��y�ߢ�V)o��{P��W�U]��J�8x��ӄ1�zZ�ݤ7{*NF��`tJY���)�@��o��8��)i͠/����x�������4��qÆ)=�O��wnyF7��r&���FK�j�QTo	��ja2��6Rǝ�Uŝ���&���r����@8�Ʒ����V�B�׷��)u���_�n���]���,вx���cm!_OfL�[��a'�3�$i���N#�G�\?1�0׃Z[^]G��B`Jv��w�x_��?L�Q&�:EUP73��4�ҬڵϹ��@���_�H<�PzR���(�:2}��li.����"���ȟW�w�����~�L��U3v�"k���=��eFk
�X��Թ��!'���i;����ן>��%� g(��e��ψ+��!'򴄱)b����/ϻ��C��`�H�v��o�2&����}��@P���~5�D�Gx�Fjh��񾵹xW�j��pR/�R�;Q]].��_.�N28.��GtD6:�^��W�3Q'�`�ADػ	w���/�O{x��e��m&��揔2o�"O�y#y��^�>H0D�� �|�|���id[i�У�Ocu�����5S��5:Dz���\���̾O�L}���<P[�S����d<�.z�VBE��N~o�j��B��~h�N�H�����p�F0�A�����_�0e��	]KF��-�-�c�
�S�����q,�D�ĚTR�����%Xc�o��5��^�uxd�nZ=��D�N�����bx�Ec>Y`�5ͧ$it��-�Ԫ��@~l��`�Ƴ-a�M�Q!�B,LZ@}s�+��o5���*����c�B�z F:�b3*���̤�D�����5ԗN\�fE0M��"^5Q��z#��T�Dy�V��s��Be��2��<t���oǻ+`2i��&�ZH�mu�Š"��C�O��+#�5v@��r�eWRc�@�\.�;�c��f����B�F���:�`���Hb�NB�b��o� ڈ�J�R4rL�� ���]�4c���1Ud��,Q�p=u��#%ǭ3,� �r�ށ*��5L�HY5��Ó��h�\{t"�����r��a4��:#�����T�k_�<��Ӡ�� ��V�r�2]��Z3s^B��n���o"�%��W�^�,2��ӫ'�_`��lTer��R����v&vp�\�G�����_%��e+�N�߭(�-m��/6����!_�5+tgK����n7�F��펴��7&!hK����1%�t2o�D����&�İ����0�p�2��C�V���P���c�*Qq"�]|�K5u��T�I 
���z=�1P�W�j$k#q�W#����_ú���
-/P��G�D!e.t������'��2��ಔ����� 8'���\b�F-�v����\��Wt~Xm�-����/��U譭�ƽ�2���m�H	��SOn��Q(RQ�{�@�"Q>��l��spʭX��bQh����3h�;�*��|��׼�ʷ	?���XZ\�>��t\H IH]7ɐ+
J:�".U%]�g�-���!���N׀��ҵՠHe���rR�j"-��a�Ʈ�V������)о��\�����"Rdw�1)����Ɇ{G��e�z���[��zy�n{��������؎���R����£:C1u�)W����}ٴ[(��|���T�k� ���D�{C�H������lRr��q-נ鎖-���%�tj?ܱ�*�vpԜ�J����K���ׁ��՝�᥿.}@�qjGFo�8� �r��/QsވqC@p�#|س�Y��~7��1dV�F�������F�Dt�F`��Uz����%2	�PY�fxb�f���Ic���ȫ������������Y�B�%*���n;�z�䮭�-���f�4���j���Ysq\��bՆ�EI��ٜ��	I�h�Z�`aF��
�J�#�L�i���ys�����=�\��QW�m�2��9:���?����&�JA��%�-��\J��gݗE�Slm�t߆K�	��*O��d'��͆���` �_�~�g�7c�D� ��l?ɩ?R�'�A]�T�TE�)#%��������Z�8A��T������3n���֤��Y�Њ�"h�z�o��6h<AT� �ɔ�	�M�������P��0�w��pU�τc?�H�����}Q�W-�j�#L} !��:A�"��:l^��
��C�����`-�A�cH���#߄�q��R]&�h0�>����<�.�r9T���~睍-{��3�i)e��ɂS�p�-���o��sR��������{^^�w�/z_H��3V��-F1�\���Fs	����|�>�a��
Z�t��-��� a�F�(5i#K�Y�H(7��O�E]\����sO-�s���vˊ�� ;��W�"�-$V�@0�y\MQe�$G�LCF����n?v�
2�i�Ri��a>O��}s)�����E���o�����5`��i�aFU��3s6���}Mkİwǌ�+��S�:� ���6r��"�=��Cp]�7H��	?6�
ɽ���4�٣K�G����.vP��E=.)�O2QcL��3�rr�p���+�^@|8�1P(X���Et	6��a�8��#���w��Rp��	`�	�~��^��@[��@$�7{c�F�b������^��A�T]a:y�3��x��
�n_珚r������HZ��¢|}�L'ej��@e��)�5[M"�dz�خ�`"��:�K�91��3�3�W.����C!�d�,�e�t��?〩�Om[�~|��!t�Z�>�����;�� �#Zk�m�h�����i`�nj��;��LcP02���,^�C9&nݘ@���
� M��m���^*l�#��>���±t�PW��nw��E��v�4^�~K���+�v���B������*TXV6]���I�j@qZ�2��(ܹ�u��s��U}p	��j��Wܓ���9-Y��6wz|K�
f��S�TU�����9��09�~N���`�9���<j���wD�om�\ ^�qI���6�C��w�^�%�HJ�?:��Xse� gN9���\�a�	M����vv�-�ߴ�La4_�*��tF㦥���S��BӒ½�Ԃ����I�A��ի������^$"�MY�k�l?GS���9�:��{��D���'�ryu~kjCQCNL�[�O��Ժ���T$�K �^��5�;�l�⼼;��c���]*���v�B�?M#<N�}~�e�/ڶ#o�\����f�(u�H� >�8P�T_�a��)L����)�
iM8"�ؐ����Q-�$̢E$�s�i���u������F���dh͜�_�\-c%}X,��ݛHy[k��a�^��VA\�ux$ ���C�9|r:�O��|�
�K���2���C����z���X��;����<�S2*y����~����
�A�6 ��뭤C�LP��]Q�'�]`k��pUկ܎���"���"%\9֭6��YC�߸m�@�������3����� ������B�l�J�6��`6Ϻ����稜�?�f}j�Jm�T<~�K��4)�{ ��mJ8D�SF-���i�i?^�N�H���2���G���:�<�[�N<h�R���|+��;��;���p?r���7 77�h�v��_�DMr�
�k��Ĳ��0{�aL�c�k�r���r��y�ø!�SN�D� % �(*�N�_�e�� ��lϫ#�U�!��\��VC[	�30��68������Ɵިl`�[m4"�x�43#�djG�����Pw�E�0�Z�ú�S�)յ�!?P��<���� ���k�G�_hk��	�L��<�G0y��jԵ�6%	_�q�:��ѣS�Q�~�Xl�Y�<��"�W8[­�+�b���K�!$6�����pY��Z5*�+B�_[�����	��O����5�s�FX.��B��|^��E$�=#��<� g��b]�N���ǜ�]-�J��<\�TB0Oʹ	!�%�T*�U�p�"�Btm�zó���!��.�z�����ld��W� �^$�7]I/��yڋgZAX�%M���w��uA�lKݢ����A�������4s�y�V�rUJ�\�6��%,i���_BO�{W�����<��=��n}~��X{k�՘��{��0��FU��4�nH�Cd�����2^|�]��k���oT���|�e��p���F%�,�b+NmFg҅�'��|����!��S�A��NY�q�7]�����<�Q��_^���� T���q�V�b5p�MU!O�+*��"����k6gqI��CIe�n�vn"�YW��p�2�ƫPbwUߧO�$���_0�m��cʞœSq�at@%��n���ٙ��[8C������,ZD��A[��㭷��,�R@`���>��p�����!&�r�pn�=&����+c@���g�녔ܨkX�� Ǩ+�w��+�sP�I���L߈@C����H��1����Z���<���5���9+.D����PL��Z��֬ļ�l�0"Ư�-V%o�t���P�wUV�GM�O�|m�LuT�>������fG�?}��AЕ���-��AL��Q�pv�R�~�>EXk�~��~H�ؔu�����3�+��})�ȧ��ϲ�4����A��DYĩ^)x��I�?�I��(zM_3�;gR�v���pyQ=H~O������G�Ȟ�����[}�I�'�����|�WخI�a?��Tn�ŏ����}%��#�>0O�Ӫ+o������#�!M1~�.�����E��Z0L�A��g�§�0��	��vv�/]�"��>��o��j0τyu�knO��Ɩ�J
vzn����ެ�����d9^9aY%+i�j�`�T�6Ɓd
����s+�q������'�W̮IE')��Л��K/�����9knT�zo�Hr:�ɎԟX��O���`&�o8����.�Vֽ0� t��iˏ�� _�m�&\�Kk )���q(](O"�1ŗJ�TM{�)�G�oNk���[��Or�	9퀻q�{��Y4����<�����kbG&����I�
(\טC�^N.�d�593!0ߍ��r��<��p"o��y~�L��<_��)�&��WO,�3���@M����h���T�Ɠ�8��t��b1�CYU�О�^O��[B}t3F~\V���N<��0����֦:h�i3	��S����v��0hz�����j�}�+��|��>����4������NcO��8���'�.K�PVk��+z͏�w�%�6F#]W��\�J���ȴ��]6��j�m,hn-B+�n�	�	w�[$@n��j)y�[�w�]���s'�dكN\4_,��J3$'߂���	D�z�6�����^���p5\6;3��P޿�h���g�:�3�����MJ9���B`���Xkq�XY��o���~���w�����őDw{H~��9h���r�1�}��#��;x��߮2v�cX��Ά"��t�O���3�,nD�iƌ��D�dSN0A�Q�&b,��1Zgi�;���I�sw"o � �f ���yo�"	��e��%��"M�86��Ν|��ӿ����.�{YI�W��qK��H�AӃf�&>�8j(.��������.�i\<�pRe����5���Ϸ�Ӥ�O?��d7�ϜoK��I�p�Xl��7 ���?�)Q�a!ǿ~�4)�o"i��m��� ����lLZ����)s�\_�����v�����M���4���A	��
���xC8e˰7�A�h���'�ߟ�u �����4��ka�Nf��k�.xm`�j�&=�)_g4�~V���n�c]�;n;�X����N:����ˑ� 5ŝ��~n�p4�,�x�-�3V���ՃUpr��h�H{JN�Y�!`(@c�>᰸��s�՜�=� ���;��zp�z����ۃX�R#��)|��qul��-tHG�{Xb�h9!���.~N�1Pf��J��E:[I�5x�0✉N޸|ms�D�Ώ�Ǝ�L|6�W��	��� �sA�\&@�M8CQsFu�& _�#J�S��Z�
�����8^_�:G�H)g�VU��\�<&���r��m��4H�����HU�s`$`�&ں�lƆ�͝�o$b!��D>$����yP��v�Z%��%,��Z���JT���,<�-�;:��c�L��h
a^�~�㰱�e;�+���@d�o��O�?���߳�E�þ�U���/��vO��;�D%��E�]���w��� e�>A���)��+-��sSv�Zݿ�+5�Qּ�hgd�N�%ƌ9��#1	���1w��$�ݒ���N�Z��Qg��	R������q���Y���ro�|吀��&�y���֬�0��X&^bDܿ�p{F��wA�쩑�i�u�����ԿDg�G'�1�I��4f�X����Ul��������>M�Ms��B>�9ua���^3ߺ�	�4=��Is����m���R�A��]��"��;����3(����"��O_��~�{A�$���z��x�e�7�������z����x�-�FU9M�BGQ�_����x�ii�:�"�[�-����&'�+�@��!}�v.���O���d�%}��[�tBxX,r�S��
@6U���!�B��io1��֧�l{\���Ty����	��_�xT0�v[�{�{4�8�ؖ����:D؞ua;ѹ�ݩ�.���r���W�_�WY2��tgoL�u>K��WKϾ���^-��P� ̀_�)v�-�,>�4x�ƭ.��eŶ�.��v���&X��=J��&B�!�H'f&ŕ9 H�_!tV��2{�\l����h�3Q@[τ*]7�
�����$�}_>:�"#ө:K��9�N�J=��y�7�@���7"Rm���)#�ЙL����E\=/ZĞ��2Ċ�� pv*
�/�9���[�k��+m���O��.()�����]�	-@-B��*��3 ��	����d�4M�N� 4n������8a�������F`���CTSRc}��bQbBKQҧ�&�VݙID	�[}Mk&�2�o'D��Я6�u��� Fpq-,,��H���Ђ'&6�����2�(��>����u���0���t���)�� �`���~R�%�qEc}�&�6Z�P7x<�_J�<�K��w+k�ӓ����W���Pe��l3\��3��\�؆%C� �f�e/ț�������[,!�2���n��^��_�?�t9m�(�BeW/2�C�2����F��i[vS#�@,o1�{���z�36\$��fV��-^>QU���dV���\�U���+�\�C�!����Ͽ���O�9^�~�j	"�ӭ�0E5w��ܦ�Q�Jt�q ��:�9Չ˭;w= �7'h�:�e
o_����~za��9�n��z�u��o��iNh�f�s4b�7�˪�jEF�w1��t>3�5��Hע�;�/V��M��S�]�Iu�C9p&�{��2��r�?/�6-����~���V��Q��T���g���r�\�}R6��5Z���ah#�C��o��'�x*yA߸&XlxV64EB    567f     8f0�O-ӭ#�U�:��`���x`;V�I������:�v�X��|� G�D��P�DGA�e���,�j�.�ć����	Y:�3�Q�1A��Q��ŗj�������q׉�ܽ�����KF~E��Uc�.`ǧ�nuͺ�Vw�0�G�4��/>úE bk�=̕G�ƿ�dU:}b�U�)(n�?��++/��]���5�8�t�Д�G��Аg�*|�.3�'e�K����|��!�M�/�q^ٻ�lR&k��X,IyD����Y��ص)���Q"v�},92�5P\c�������ܬH�ʬo�e����m*� C�!"���;7�����cZ��F#�ͣ�]��%y��X2X���W��F1^�G�ˠ\CWH�'�|6U����P��ܡ��.a�wH�s������Y49`�H�F�O7Y���eJ@�F�kz���$}>�@19L�-C�M�m�Awg�ߵyP���]�� >Z�E��5�Y��7�<\T1������iQC3���>und�Q;G�	�̩��@+a�?X��J�IE��0������0�H����J�7, 92�S�vz�����Ś ��<�2[Ϝ�o��q惝�zy'����
+���$fϚp����􅔘���:�����%�ڸ����b�{jk= �+���?���CViqQ-[Y�_/��P��YT�kY1_��ۭ"<L	,m�IDg��uҤ"�dȆ�8�B|�-��&�XI+���j�������>�_HD�6���1)��ަ4��%�e��<yy���Ώ���R9�>�4�u�a�O���(���{���
��`���mm~�0ajR��K��h���5����Fs�	���4e�e�y�{��\�; ��ܪ��FL )�dQ�Ng<9�'qk��"���p4����%dOID�/�tWN��%*�po$0LB�z�8�)U�|�WK!\�Y�T.�N�V��v,ޢط�D�i��dy`�� ����y=�� E�������P��+��f 	�!�����C� 'Щq��|�E�j����'}U���b9R��{�>�l�J_t��)�H�N�j�˷:zB���r��#�l���"i}ȹ1�~2X@worT;y�P"�ck;;b�P�2����v���$�~�C��U8�kXv�ɴ�.C~����x���I��ѪҹrmX���?��}�Ɠ�sa�b����s����$�����4%��x5\a��/1w|��p~�$�3�7��Hm�+ӟ\?�L�>�	�f����9���8��!2���36HHi��՟5�CB�5*�D"�@��9��n�-�2���W�{�	�ʝ2���h�� ��T"9��2U<%@$�`Mͽ�� ��g-3������	Db�s�d79�e,9櫕hX#�`�K[ 'P�	hS�L7��"�p�)�/�G�wl�s��N�� ��Y������S�2�L��a�x��߲{��eŏ�١�Tv8-Sdt�zy���>Y�s��z�O[��0fl��GZB_rk�ORO��c[�����Hq2��E_�)M�mƨ��ҽ}=�x�欁?��6ċ����1?--�T;�<����p{pN��\)V�kv?eM�z����;ۉb �1A�J	�C��/Χ*X�JGxva�?�#A-(��|Ѽܧ1Y)���8���6�����b����� ԏ��X�� ����֬�@C�#�5��q7S-9�:R�~�mL����t�V�iJ'l%	�83���x�����UԌb9��ͳ���KR*��av��gOU�!��!��H�<�����b4��X{�ؤ�f|ЇK�D[-����[pSC)��Lb����u{�ʉ?��'��Č���VT2�O�|�D�����|���2Do��"/=�xΖw��&(گDG�	���\ӫ(� �8A-�Woa�6b�re���t����_�h�����o�A)�ψ���ݸ�]#2�&�]1Sw�5��
�G�����Û]ad$t������+�6�F�k��4��ς2`vE7�#~yMxy���8 w֬�I f���5e�x,�{��o��7��1�������z��Z?
��ʵ:��D�p/��!-��g������ &�2?�[j��nJO��\��/��k�*��m�s�6�,���ӣ�a5=X�Y�=I�*��1���ku��t�����)��տ�b�1���R�6�#�����RZ�wR{vʍ�>̦?���h����!]u����K({;|�?����˾L����