XlxV64EB    1727     870�̞g�Q�MlP�w!o���0u���4���=���جh���!����[�,`�p9������=H4�5{�M�
�,�<N g%��� �7/�B�}8��(#��J�<yU����g��ۊu�w���}���b�E��xkf[,�{���y�1N8�qbŴ܏�cM/^o���Gr�Z���O��@�7��4i�f0G?��k$F �L#��������o�a�[ì���G�B\�^�����/�y���c�$�~,�'a7H���M�}�@T�D�w���|��t���f���Γ�Ǩ������*VdBF ����5���b:�,��SWx0�C��ت�E`�j�]�\	��bsW3�ߦ3�]�L�N�+��A����� �_5��3�a<VX��!#�Y�w��޼�m��� �7��V�L��F���J�f0��u 9^e����>&pY�'w]�w�����NPyII�]
� ��,�tε�P����vz�7$��Q�^u�DO�>�cݳ4j^��&8$�9�Hw*{��8���$r���J4[�=����M��j�V^Y��f����xf��*�! ��!��˓�Q�#T zxN�P��4eU0fw_)��w��Y_.�o�W�x^�r`���vrq�{��L�%����뼏8�b������A2<%���uwJ�?�C�+����I�z��~��Z��"�X%���Nʃ���{���|�rzԘҒ����@?4f�2z����v�C�:��5��*�����~L��)���2&B��)�`�wi���a��F�)��н@�k���'�\��>K��e�N��"�.U������_d+D(�"����tk����t_p�l��/Θ5$����j�A�/�^�d�^�mrֈ���MN��v|W.͜�e�
��s���g�x�y�8��hy�p�8��?���ٸ�����
۞ۥ�1�S�q�0�6dd*su�Z�Jb�7�w���ڥŔjg��>�M���j���k8���9.Z�s���GO���rm�}$<�7k�\$��eEOa7��*�1���Q����?^��r�s�pQ��i��\�>�݀ǽ�m*�qE� zMEu3��V������Ł��l��"��R�H�g�O�2�KRް=�ԒH�Wi����I��k
��e�4tEv�-��_+ڇo�J�ey���2�x��XL ���`�T�&�35����c����ci�3����k�0�y�/2�T_���L}l:`�⵱���ڳ���įu�?lM�䱃s���B�g[ɝ	~\��XP8�����-R]����D��"��m��e ���A�.7v��v�2l ���2J�ʘ��N�n��o�t�H%�G���
�s�kVl��Oj��$���<A��#�O�tM(%)��^H9O?�/��cF������jr��ӧ>��~򸀒���nΰ��4L\Ēr�:��8���Ӻ[~X갾s�.����ܠZ��L����{9���{[o�]�R��'���p�0tSڧ:����ȝ���2h4�����?��%df���D�xj��GR]%R<�W�t`�O΄��~��.��`9��Z�+�Y���U�5]�$�	��ی^�����Y�H��{�Y/ؕ��֛wVh�q�������.r�x���Kk��$6��aZ� ��G-⩍�-9a'
��epaOU��b�y{Ȏ�W'��"Odq(w%�w��&ʟF�8{�����pgqgU������u��$�a��?�Ɨ�O���n����b�@$�HS��9�b�M$L8�n�	D+�z���Id���k(E���hc����$rԔND}$J�	�F=� � �K�=�v���G�wwQ8�)�!z���]~WZ���oH����Z�݇����:a	>�yKS�}�(ʙ)�KʭM�� �-#�|�\������՝����	м?E���.�Z`8��v���i��A�Q���
��-?�A}�Ŕ�u��5������p�+%Pc��`� �-�jR���-Ǐ.t����Rx�@2�7�'�������O݇��s� � �{��n���M�A����}gЂ���p4é�����i��G�u��i��Er!�g����.D�Ũ�ӱ��6�;���l���P*֌S��