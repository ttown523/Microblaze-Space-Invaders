XlxV64EB    1f78     9e0�a��6��aJ��T��	z3PI��֑1À��2R;�t�Z�n�r�'�;����U�yL�{�M@Z#i�x�E�8v7A��RT�42Y!��I&eՓ�
>�G��M�y�7ѽ��{�Y`q:lL��?p��̭���{ ��s��x2���9�ثD�f~:����A�����U[c�go�#�nmS�TT(����nG����/�rbd^i��><>�V4�m�=��~4�����0sǙm���� ��D�lM�`q�pʝy�*?��k��S^���e9s�E���	Șע�00It�},�v%�76�<�3��!j���-�F�4������/��{�6���I���J���X�x�p0!}�J8ş�LE�/<׫�lהީ
�tk�zEY&�]��e��gQ�=fyF~�kցk8��t�,�}}��t;�oő�B���▦I���e�Ӑ6����_�N��7�ˇ�C�}!�9gy�R,đ�V�h���⵮��'����ſ=���+%.Ť6ٯ^1���h�1���LG36\���N�f+k�+"�}U�eY�F|�n��h�0LY}���H�~��D���o700��gT�9,�#��6^&�G9Iη�y<
C,��\a��o�L����j���;Tj(�jCw
� C�0I�A/7�����&by=>�|Y�y}�`�@>,	��Y~��
��َA�5d��S�6����/��н�e֝�e���W`�!q�AqB۔��g���w�C����<�GѕI�go�Y�~��y��WDCE�1��	BB��Z�^8��Fq�Q��jw�grZ
@��Z5��6�H[��6����<�~Y'k�!T-�K��4Z TC�ZQ8�F|�*�n��75w����"`��3l'_$�q�0P���A]�AVj�&M6��\_0�@�2?$Q�qK���{|�)l���{�_�~�"8�5.[���@�ʃp%N������6 ��
a�SH�-4��Q�� #q�L,���A��; �I�Ď�K�g�
c��������Ū覤�Ä߫� ޯh�*69�Z�}�t�t��p����1��6��pF���娛��pJ��Z��y7�3������D�(4��!��h����DEn̙�l�~>uRm���x絭��z�U8J�j�oN��0=�1���H/��E����>�'�W��.�B\`8H׬P?
Z�#��xj�FUL�dNe5����������PodX���鎌�g#�麳���G��'���=��"a���M�������3�W�?�(YF1ͱR;�G��$!�Ě�Z_6S��s�/h�,�t4�O��e|�.-G#F4gr��
�:w�FV%ƻ3�>�i�E@��	��p�:�(D��9�?r%��n���P��@���P�7�)ڽ�Nw���~ÒWX�V1�l9�"���Gmw������/�8��*�m����-�ٕ�A�G�jE2��R����ɹTP* �x��=u��6��鬔r��c�8�ӆ��݌vb�xe7ap�XáA���x��� �n}v�r&�;��&���7fL~;m�`�壃�%<\�m�K--̭��ł�m ��F�)$4+�	��I��vy.�% w�cs���Ņ�'N�h{B��A����p�D�9�d�b�l
f�1�|�ɫ�G�hLdT_��>���ۏ���$X�",%.��Ό��7,
AP�]�R*��Z��M C8zP`ԕ��י���"h�*;]���
�NiiOB���sN�Y�C�(�͔�W�ԴG�s�����Z{8;;�/O���n��D:�f���O���XI�V�g�܋�����n0����st.��3�e衴�k��l(/��#����w<nO�}�r񮖞������x�����I2�S?\�@"Ak�G�M]�5KG�#�H5̲`7?ߡ�w�db�t)��b����D#�� �����U�ȉ�|�_��S.\B-rԛ/�H<8�8z���
b��N���3���)rf���{�%��@pڍ�?�r�$�ʪ-}���\��	��P6�����������^���N9��ͮ�қ'�ٯ�J��G=ĉ)�~����^��8/�Zg��o���vwhj���Yvp�����H���`.�ʗQ���"3� ��
K���@�N㖢��¶$�����d,�v ݺ�:ψo���,��?~�̮�8 R�t�=��sa��,�����KO2_��/GȀ��C�\�T��r�K��Z$5�H���	�&a9�]-���D�|������Q�����0^Ѡ��8@1⏴��S9L���d�ԇѶ*�}%5s���}�'���D�Ww��{�����g��GZ����)�ʾ���A�ld	ĥ���J���K��$
�g{��]w�@Z�M��b��:f����%����<	8e���	�Od��q��k-�=��>���xm�#Md斠�]Z�\s�W��Z����L�u 0X�K��f��>V����'�n~���(;�WL