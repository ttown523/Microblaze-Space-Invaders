XlxV64EB    1b83     9c05��R�=H���@���:���9`�=	�hzqb�����	Y�hf�T����Ym�=�ճ>�\��>5jB�F�g3(I��+h�Z3u	��:�E��̗6�s �Tf��YmZ>�td�v���ѵ������|f/�>~����y���$����A[sSWَԗOc�w%3����Gf��7\=��"���E�@�]kGE�b;ӈ���0�oF�9c��|L=�����m�Q*Va�>����&5ZC�x�)絸@<� ���Ab����`��#�N�DZבs��S��� �V���$� �g���n�eYC	ߖgo�>㉌��#UW�������v�]��)U&��3��Z����.�(�QPm��ғ��v�2�`�{����q��;oپ���Q��u�n�j�����8 ���J���nY� ��bYh��s���	&A���N`��n�T��!�&ȃ�C�[���S��p�aY6��Zg:LѵUxT��Y�� ��*���T�_��ʤ��v�K�Z�8�jo��� :_��3A� �W�kp���+	�j�\p� |������'˗���
��^k�m-�Q�.�we!;�@V&�U<`|��|��s�G-E˶��i����j��d�T�QÒl��ﮋC�_E�u.�z�\Y����p�R�7�+��iJ+b͇4�e"�U��F�*9'�F�5�赼l�5�M
��n��SJ̎;}�<%j�h~$��j$���p�H+������e�C���1��n��EpsC�q��r"&����X �2��H�x`��Ś���;�������)je=`����eϴu���h�llޥP"1X�`c��`^U�&�B���QnF��w��H���kO/���9�A�D����6	��q7�NG\6ϧ�m�v��x{5-�$	^��
�?s��{c�J!�H�yͲo�� ����V��cW��7�O��Rd��],��M��.�p�_c�gc�+�mQ����
-{P�3C�B��IhL~"k��Z�o�d�)�G��'�v�[���j�6�咖�e�$U�j%5Ĳ3,����[8��3��+���Rz�E�Z#FS+NEݤEB��m�o�6z|�ڃ�	C:��փn_���8�q��	ƕo�:��@\�P�Ab�n?d�k{g�]��52V�@S�1�0uDU+�	pV[�l��t�$�0����G�Ak����$�9������B���� ��hKA���=�_�ߦ��cy٫ƃ٨X��kPE�#�Խ-:)q���5���@ 04$1;`��7�T2������-��Z�D��.�-HW)�)�ƣ��_���JX��!D�R�m�p��cA*t��b���G�P������M�3�A&o՟��n���&�ճ�`5F:�a]b�Hz�V����5{�^�n��ċ���	�FN�g��G����+��q4["�Ӝ�m�9� �X����8Bׯ�C�CvI�[BDu.dxj1l�}��Oz������G��Z��h�݉��z�z��������a��i���zs���q �4��yC	�%P�O����١i	o��V��nAp�C��_��,�"�GS5�>�����k�nĝl������{H&v�Px��{����./��+p��L����t9cF�VbK�1���e�|�䝪���U�I�h|�{t�#3o	>-Ų�6�!S:�a)Qt�e?�HOχ�sZ���6|�5���W��zw	)�m/R&��(����o����Ni^�{s31l�>4����O�^��۪q�Z,ʿ�[{bj�x4��9010���F�����=��L]
�NW.���8_�]֯?n��M��������G��|q�I���%xW��QVJ���7����,���}�bxi�p8��a�0����i�:��	�Dd�����
����piU����.X�Ґ���cA+hC)g�}�ͺZ��:ɛ�]|`Spr����#~�Q[/X����Am�s.۩�u}�`�^�)�r�+�y��ܔٮ��{L	����SR�8�u�e3�	��K�[�K��Rzm��'h �0���屠�o�������'�'in��B1a�S,c������*h��!<�`��>V%䯨�[J�0�����a?_��m��s��h��Aӕ�C�[z�	!��a��M�&h�Z��Yw��P��HPc���f}��[K���މm�#�9����;��KS_/��4_*�\��#�C�m8�_���r��*�L���<�����o�Vn� (IY�c����g�Fn�~�#��n���(ϵ<4mn����z��(!爜/�z��<��y҅����&��`e�e���JS�-���
k��#��f%��c3	d���m�R�^���ݹ�<�i�93Aּ�*mQ,ĺl3�W�ߋ�D߆�30"imv��ċO�ey�7�2'|����H1<Г95�X��y[��