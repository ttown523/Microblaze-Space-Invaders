XlxV64EB    5dc3    1420��������?a`TX��<K�H&v����a�& C�[~��Ϧ>���Ӯ*2�_�{t�(�����6H�8`)\�v����{��#��):�l�KR<��	�.s�|kԊ�䐟~��(\h46�@�MOϒ�5<B�g�I��S[a���
�seip�1�с�����1(�qQh~)�Ù*����l%e���\J_d��Ґ��F
��Q�5����cZ��4\�eQ���5��K��n�F,�~���K��'?]ٕ�YQ�}?���xnںR�_휚�d�gI��< Xd��Y�B���DzE}0Fj�<�%�I;��'	�g@b?[QӯW�kc�m��`��=�KD��t���݉�G ���%�}�¼�42��Ѻ�����W��		A��w@}�y_@�j��D��)����j:��]�fA�tx��g��a���̷����v�ĳ�l2I�}�$D��Z;�6\�l��ie�4(�_� �`�`	��K+�o�p���x$H�w�@�	��n�A]�в��oW1�}��G/Fw��^�h�v�:�S���i���F�^��6�����=C�m#�*�3����Iulmy䵎�[o;O�4!˴��h��`��/q~._�fڈ_�8��h?@3��y��&�w^t6�o�j�^���}��E>��(Y�^ŭg��9������I�,}��9��Pt�P[ʊ:�W�[��Pr�_�rJ�@�T(�kS{>K��a�*��=o���뼿�ɆVဘP0B�eI�����/ ���hl���>@�,��q��q���R�vuEY�'O�m�2�1�Hf��$��܁��,��w�*�(���}`0�Qc*��=�!��1S����H�߳�f�MzQ�6�^a��)\�>��o�w��y��ǇC�Jߚ�������D�%pu��{��ߵx�'�yY�@~�!���~A�)[%�:̏�ѳ����U����?S;qe��W������X=����D���N���NN!���	S|j���8	ZI@ȩ��IR���hι��0�{��>���FG��igL+>��I����XR��=�����#n�o*�?MH[�_;)f���mD�.��x�il����+�,�ܙ�櫟����v�	��|��K��/��^ۗG�c�I�\�n�r�b�5=-f{��6�rE�CJ�H{{���Ӯf��:l �7��Y/\xȹ�棲�B((�.�]!**��+�"2#���<�5�uc\SA���C"����z1K�z�v<����HD2�k����Q%UX�'�-���,�{�H���|r��O�}b���O�1�v�bA]�j���
̆��ݙ�>��^M
��#�9\{�;k�!� ���׼���b�h�d�s	h�/�c]j�G����Z��p�����:H�P�|I4d�����ܓ�Dl����=��@�~��^�����*����������Ǆ����Z��W�-z�`�U��l��g�j%�����ݻΛ���1�0�v��n�G�f�7ij�bRB�`>��|�
/����J׿����V��N(�H��KM?�!emaY]��Z�b���?j���'l��
����ݴ"�?�]`�Jvx=�gǊ��Hk[���g��$�� �$ZN뼙vd�U{C���O�&\%�On��͜(�{�Cd�O>cl?�TB���k;lH���a b*���QK��I#��$�������.�4���c'��/�&�Ap�G�T��g�r�b9O*�[ v�2�Lb�t{O'Q �iœ�ՠ]PԪ2��Ry���E�0��6U��7���q�,숯�,��~�����aL:���ty
�����Q��Ci�/ަ6َ��?�ٚ������d!A�j�dW�B�QG�ݰ�VA�Ug��l�ѩ�y�i*���؈�f�S�����廉�p����m�����,�3���V=ƙ1�-O4��.�嫥p��:�`f�yE�:.�qq�S{�O6ek�n����d�R��Ҏ�M�zT��u,	�+rnp=̓�Hb�{>A�8v����7�1�(�n�Lf�7ϳ��A�*�K�~Tb��Ŵά��Ўֻ�ϣ:�W��\�����
��{(E	N�;�d�BU�̊!��K�H�7�n�'74�&�(at9υ��z�ܹ���q��~om�[��_f��o�,>0��@����W?�g�%`&�cb��\�򓑠�w�1���D>�E$�`��Y�F��U�4Q��l��������믟�Q�kb���k����}go�%R��=t=5t����F&�.��k,K{��C�cZ+Ѕx ��tK��<Y�b���lqh�Y&\F�E�b�s�ŖfS���9G�ɘ�-��|���@�\���"����S-���x�X��C���2rܸ�i}[X/3z	��7�룧�c�T���tLz�'?8���T$��}s��X��?>�J��`�X��Ӭ��Q�5����8�f7��tC�X+�׍�u�)qc�m����[I�V�d�$�-���.��5����
m*�D?��P��q/Ou<)��ۻkt�C�m互[�m���ނ�F�V9��3�z�Η��N�D_���� ���M1����q�O�s-�|N�!q	�&� |���~�����A���lk�䰑��!l���C:ʄf)�ȉ���a��"��[o[��h_���؇���ʁ�dѵq5厢f�V��g��ph�Q���a\?����T.�ܝ�w�8�U���\�
���)�<����Nj3�X� ���
�#h��ȿ�a��m�Ř��)�W�`��P�z�"-UQn;��f0�l,8ُ�����II������؆D�*O.!8�7����Ӳ����� �*���r�f��� X ����!�A8aOo.�3��c�!'N)�J��[������Vk���~;��H�!R���^3�\�� �O�C��\fnFOkA���8�jTD���6[?���������bJ�:�xX���[j�5tF�,wX�Ǳ����[C�����߾�ޘ�0��J���V�!l��-�0�"y,«|�a��
J��[�ih�jI�m��v�9Zu)�y�&k1�{*b��s��F�`\� 8~���d�.�ӻ6�Q4�u�ߦ��7wF��2�B���^��x��}E�i�h�P��g��T,�6���U���>�1{?M�Y�=����E�Y{K-w��I��0��GB�`j���V�+��=;��؏�4i���N��VgF�=�^ �◻,���N#��淪��;��2�����f|D.���w-�%�ʕ�6��-=*	h����Ý� �b��z6�&�r�%���ׄ�Cv��%����rcVmD��R��Z�KoZ�	���RH�����ZJen��
*F	�ߜ1<#Ji@%IPWu�y�= �5~���<�s87=0/�퍽��b\]��V�{����ܣ��B���6s]w�'8�~a���lXd/�F�Χ<�vBH��oE=Oq�B�P_G�8^��j5c�"�ir� ���Х��y�%u�����X��&r��(�������l����Ĝt�+o�~�=��胵��XV�
'l��*�B�	?��0�����R��^ �ؗ����H'wɜ]�Q`Dwd-�_�6z7�zn1n7e��~�=W�Y^iM@���fሞQ[��6�c���AF���0b�M�e
��!�3�A�FU:4Q��!h"�/'�T���|?.*gܢA]a���NK$^�Q�����R��w7b��H�S��R���J{71w氌����.:��{'9i��o�#9T�v�� �X�'��b��;K!8a�&�ġw$�=<�3B�"}�_�tX��U��߹hk��( ��,��s��ͿE����$藳�!i�]���~���!ɼ����S�3P3�b덣b����Fb}
/U¡����2:<��$q,CX���	�b��|8v�RO8h�}��*�0��A��� ��=�3�Jh��pZE��&e�
�B����`�C P�p���/s�3DT��[�A��%}�C�ū�r� �-����H���UlE�Q;�!�H,�D��Q9�f�59d�¬Dy�i:�c�T|k���+p��B��d�	
]��2�k���'����&�h�vª��{ÂV���ry������P��]�̕,>�<�v��j�i�}m<�b7�e��f��_�ڤ
��Q��q&WRQ�����׊U�2��ƊGx����Sٌ��q���9��nG�9{�/�Ck��|�9�N���ی�l#N�`ƶ���>Ǝ'9u���{��y�":���9��,�w�PD�ǻ���|zKN#���;b�7S���NGGJT1~�R՜�[�"�_C)�`l��b顷���Xܿ�~:�i'���|���أ?z��-��w�T���X�8K�� �R��u!����ZA�G�wO�L�=[�};�+nͧ9��x�-�z�na4D��_�Kso��&��a	_��}CL�W�'�����h�8�����7)��tρ47�$q���oO�Xv3���H	a[��a��'��[�~�����Uz��W��	��
�����eF���d6�j���Q��#\S�:K����̬��6\���R����cex�»,}F���ZN;�:#�n�W��a�F{���Dn�6���̚�q1p2����s����u��I�ې��:�6�}w,�B��|��.���>�2�y�""ȃ0��N!$��� +��Xt�	�JD$�E-����Cz��=!թ8�
6k���Z�7Fth3g[�Хm��:6yy�ɇo�~��=�JJ�jÕ�۪�v߈J�����s�,<h'c�Ax�oO�f�=لǨq����"��	�5���{""~��=�ZH�D���Les�z�W�0���z4����w���t�Tb�u����p˼R3�C�_b�=�Vy[DhŪY��E�e����Fj߳����1&F�J�B������g�6H���(�57�N��3i�*r�4*.%"����Wg�..���Q�"��ǥ