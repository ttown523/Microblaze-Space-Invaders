XlxV64EB    2965     c00���4�A�� � ��?����t�s���p ��>(R�`�'��x�"�)�U��e^��v:�>Y��D)���\����:I�u��T�G���6���r=��]�SК�k���Q,����Ii������y��E�8'1V�k(�>(��w�a�Z��B�.�@ܳB���N��7�Vq\C���W���:�T�f��Ӏ6s�cq}�̶���M���v��9���f42�ߝD�~��O/��O��j/_�k%1�S%zz���j`�������w�V�YocAй��#���\ES��P��b��p� R��N����rm��v�%���*���|�by��}�/ad] ������/r��g���}1����Z[US%�#��+����V��Dv���̛�gQv�o� D ��aթ���$ �g�9��6`��um�6��Hƞ�c0�}�Ю�F�%�Hs��P�
뚋G��Nȃ�v�,_���U?|ӵ綁��NQE����~Ɯ�OUPi4L�6>��A���6��&�������Y?��ݝ�c0�\Js!�o�+�J�f�j����c�`�����H�����SE���5���V��튋6���Ty���2�ye�Yf���������Dר��� T!��������p�~�ip�E�#y)�l�э���ý	k�A�P&�6�KB2�Ka�!��j�% ��g�u �G�D���s��LTǃ�g���j�\T�A���i�C�K���w�Յ|�=��<i[[ߞ��z�6�%�	��� 4�]Q�4m�P39�h��j�oEo�SKI�Q+��>Sv⨱ �-Tw��'lY��zX�x�� ��w`Ƨe�,�c�RS ����W<Þx]L|o�Pլ���v �׫�n�D�� ��@��F��D�Y��W�6=�9����>�b%�h���R�c~�y�L�N�<�;%�?��Wu.��Ҋ,��f�V�ѰL��W�_��Au'��۾� ��#���nH�^ֿ�}�,u_������|H6�� �vco[��9��ℙ�m�ف Iͨ<	N��as�?7a���6>4�f�^����%	?��*P ����?��Q���R�fA�L�p��C)V>��'a�g���� �Vtj��8�1\�/�W�]��k5;��<)܄�'����앿K�t�5�7���6�l��e0�N
�(ୖj]<kuɸ�� ��e�!�j���8�J|�
1eǊ�~�g�6�[�$f�_��wZ�*K��n>cct	O_�����,���]-RJ�b4'w#���1�AD�b.JN����<�
�i{��uw-�_r;*����3�f� ���q�<7���S�c (����>��d[��IOs|�Ɉ� y L���N�&N�6߆�.�͋�R���2i�+�f��7_�f�������ʛZ���J�\ 4��֫����9�H�T*�1r���t=#��r�� �b�i��߮���+A�������Z�/�`ق�@v��op�%/�R�w}�,2݈�W�������ߙտ�+�G�0�,9�2�%�P��t��"_M!�5dqGtt[������	�X/�Y�Q{�f�
���v� U��s��l[�K�R�4~4��}#F��?;��`�(��(N'W�j���T�.g�@�д�m~��1UJiLhj��)���G�DF�-�(����'7����0�߈w�;6ůV1�ܓ�8P����uCE�����r��>liO�ϭR��B�p��EwSr�Lҍo�3�v�������.�
��5�hl�*l��x3t�j������L�Ƶ&��z�	NE�1w�퍸��m'�BE�97�� ��r|��4]j�ٛ�DO��
���Lv�oz��%7�s�yh�F�V�"����L�gAG����यc���Ap-���q	�t�R�2���z�����T�i�D)�@D1r�(����S�ģ����������
4�_],	=?��8h�t�5\䨮��73��2�Z�.+��q�'Ej�	��M��GA��f��4U��?j��A��P��H���@T�9ٶ�6����cB�=2��δQ��>g�dh�15�3~R��g�b���3��,��N�a��"��{.F2@�[6_5G�O=.�Nk�6[�[A�`��S ֑��ZYy����˳".ċQ	BG��G�����E'�(\p����0^���?g+x����(d��N��e�7��W�o5���i�vĀ� ֲ�M�1��q���Ee=�B'��|�b�M�涮�����.��\j% k����W-��>�ӧB92��+q�sm�_���|���C��R^g���=v�<'�#i������[qe�,J��㧢a���+>Y���ql�ؚ�h=5��/�C��ñ���2�����l����^,�xgb_���������/;��V�����	��rq71�[h\,&�����u����W�9v�Q��+�)�+�)�Hcx������=�N��B���YZ���}��(U5�Ml gl���ɾO	mKp��o_��ϣw�eK�C2��BnژI�X�܌NMb}�y[�ˇ2��5l0�X�$6�o�"ˁ2P��݆AlSY:���.���9%��q�3�(z~��Y��X�%l}���%6�>�,u=a=EG �����5>�:�lt;ư7u��˟M@�}$���#�ޖ�����'u[���8��50��|��X�&�k<�5@�R"�x��UڱFL�PZ���xw[]��Q%�@�bȿ��M�Y�iӵt�����G��(�>i@� Y�s��w�U��cj��<�x[����b���)��	"ɗq�I��m$�c���sru����Q��xy�L�ozsU՞�`�3���{@j�H0�߂�<	1�n���1�a�S%-��h7T��pa:$"K���F�,U�I���Hm~%�`���n-Q�.�a��Oi�BW��x�r��L֎ɣDy�X+�0S)�+~ƞ\�R��"n�t5��j(�y8]��Ū ~�9E�F�ֺ�e�+��b�ײ3�