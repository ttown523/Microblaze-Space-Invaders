XlxV64EB    39d7     f10H�Z�jg�iܞ���X�^����N(mc$;�jY5�'�L��\~B-��m��� ���N�N�������24��\���n����4�����"����}�|a��W��'���y���l�ti_iP��+ z� W�3�Tb5aN�D�hD�E�y_-[�<̆(�$KF��j�+�soJ�e����y|ٮ�1 ���U��M�*�P�)�;���hO�KN�T{_�^W6JiG�
-�0H�|3��։<ks�"t��zK'��?Du���#o^{�^H���\2�m��gL^�y�zG����Ë�/3t]��XW�X�����)K�jo�`�'O>�鹎�vAݣRO'Xf妄K�y�tJ|^*��y������Ab�X�G�]��ऑ��>0e�'���E�)�0Y��O�f6�:�� @�,I�O���w'a�z��sGM$��L`�J����U��:$t����8���K�C�/Q�+C�e�Huj`����[1����k�Mߌ��D�d��;1��I2ei���i�v%�ok?��?����6�H�� �(���;���~p�y�}�^4���-MnB�\Q����%��*qI�G�񲃋f�]uS�y�z�cG����aI���CV���͍M��ɖݮ���x��F���h�H_��,�,��Ç�P� ��X�%4p�6�W�ld�h���X�e8C��Z����8�&�-u�-�و�	�Q�-��^p��U�D|�dj�����t@�t�G�Ӗ�ccQ���#���Q�f|@u��p�]|��C�c�k4嘔�����\�rrj��U@m�剜�{"e�7�x ���_�� ��9U�R����_�ҡ��8��Z�UO#[��Az-*Α�6>:<n��G��4l �R��M1{���c����o��#�~.�#3���o7f1U܈7�Ux�1j�'}�s��U�џ�^����L�4����c(�ǣ�v{�c��ܹ�	,�7�d�%�E�HF�=mvu����"DA�o�@y�idr�C�uL>c$$ڄ����$��g���A��/d�J�>^+J���b<z�A�����@���z3��>YB�y]y������Ec7/���H:�%�ppnB>���������iSa"�qӄ+���_�ׅ�f�un.t�����lg�5�����wN��.���dQ�F��Ȓ���Ef��2}�5�b��7.�(��z��5?�t��g˵o�\'�q�1�蔦�DRk��7_$�LL�Aޝ�͖��ݶe��rF<x;�����v~��Q��ޫ����5���X�@�Z�3��?�ڢ%���G	�H�QB��P��Y��:�Ւ�M*Cm���}�h@���q-yR�0�- ��ڳ��H�K��,Y+���N.K`����)y0�M�`�4�[aO��Ua+�I�d��Gt�>��r�fM�Rk!Jq}�-C�|�}㵫�ۥ���������𬤡,3A��n�����ͪd�oT���Y齽n� f'�R:��;Mz�OCQ��w��oL����i3�diPڃm&�DZu7�{��5�Q9��W�+�>X���8�����ceh1��û!YΫA��ŵ�L���nE�\A$yJ<�vnp�ս!4�N��Ԏ���:�'�QjL�CP嚠����ʔ�]�)%JǪ�=9����'�e:���YjF�d�w�㛈q'�$P��
�n_��ZH^�������u�`]-"^����פ�8����10�,�(TL�
��q���br�;���]|�3D�I83�X&�����c�A��h����_������b�u+�U��aS�8F��=�_����[��CsT�e�[��$�*H����Y���,C�6@��MQEm�<��#�gCy�����H���-�8���eb�������؄�!���Z������V #\���Y���M*�K�CET�ڦ��t35�WAP!"B�"��):�#��xl�m}��%��1�
t{�/���:����Hx<|���FY�XU�D�&n��%�O|�qm�T>����d0ht�u?�o��?q~ 覫e�(���@@w�875a�Z�O���6EzYa�vH��%1�^��ֿ!�#z�I��	OvaD�d���:���g�+�ΐ/Cq�s�J����3Eq��X�C���2�q��b�F�޺n������eڋuu_����,�Y����K/7�?B>�]�w� EՔ�ѿ�[��L�z�A��v(��c�yFGJrZ��
�m���3˻�q�鼢,���RG�5�r�F��Z�A��`P3')#o�:;����]t�/w�tD�_�5�A�N�|�ƿ�NӔ"�׏9�c�:���݃/{���e���~Fոa�����Z��$��iڝ�>�ZzN�n�bh.���C���I�F���n�$���|�s;����U 
��n�c'�f���_�)�=��K�:\�"�K,��dEW����0M�O���7̯��o�<��+¶��-�vVzua�]�泑�����oY�x���B�j|�b�H����>p��I��H�n �l[���hF��:�oq4�I����#��#�"�8)�'�[�����S�@Z�S���j�.�Λ�Z�Ad�@�?Q�B#�@�Ϸ��y9cWO1RN G���}�;�pU��W��.��D"��P�\@���e&2ٚ���ǄLS�����{�K]�~�RPo/��V`���!(��!��pŵ�x|E7y��� T$ܵL��ň;��_��^���Kڥ�=?8�e�����[B���� �l����AQ�Y(�0��jwa��hT.�ʩ�_H��^L��Kٛ��!�lai���
}�>��\l"�o_;���ٓ�g��W�W�~sX���H�\|��ͬ��P�i�����������yv�%��g����V�� ���p���k�S�œs���@�uӮr�Ϭ7s�]K�i�Nf�{�V������E���v x�����4	��{��K��P��"d�D4���Y��rr��s��;]� �[�6�J��!J0m52L�S��@��s�{��$�%ʥ�U/l�A�=�AVj��?⍄�ă���`n���>�KEP���AcD�������o��`٧�M>Ez���w�X��� (�e��9L�/=�bȀ��w�0Ta���q��>���1*s4��\�gȈM��p?X�d�3�U�X��R�k=,�WQ`��j���!L��O��Vb(1�]���S�7�8"���q+z��>��E�x3�d�����@��ӊ �v9�"V,)P�(�gq��T[w��;�����/ѧ����\N�qn#�@eٸh�	�<���`��DƎE^"�U=N.y)���%Ԃw��g�f���~�x��u����%@:s����T��~�����@5��	��Gx��ݩ� �P�Q���-�],�2����E��~�˖V�B�����4���D)��� �_"��IHJAU�z�V>nK�yᵧ-�X�Y��zF�� �N���`�M�Fh��z �}�ä�E��w����i������A���f}8�`���z��X�?[p�^�2�����š�#���.�c�S7�n�v��I�z�p�s)�zV���Mj8�֨���6~M2��w���u's,4��=�_������!n�a�[�i�V��4�d����*��U��u����o�/���Ǔ	y��
���F����v�ӷN�$"ق,	4d��K��Y�o�����]p���A߱�&�\�`B�才�B�Կi[�V/����