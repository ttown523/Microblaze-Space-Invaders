XlxV64EB    3820     fc0[�V�3�3LO.��l���%AZ�`���mmB�OOf���LX2�٢㉦�6�'�e�^#%���|�{Cn��0
��� ��:���]��ࢫ-t��������� ����LP���u�/OW���M���,p	�-��>|�>7C�� �֢feB����ݢ����z��a)�����p���2��J��Q��y�DI&��n��/6���xAI�xnQ�Y���v��r]ga _�x�<�ւDo��5�k4C�]f՚5[������*�[E��D���	ktl�'����7g�����;w-�*���59���jo�r�l�&��,�yEMݱ'Y��9-vAD�\ �BI>U�X�5Z3:�2�Sq�Pk��e=֘�`�[9� B���f�9x��޷d��6�=�)r~�!'%��Ν.f��=;��ЪxRf�y��n��v���j��׼(�lB"xq��=�~^jV��'�����9�����w*y��据j\}����Wf�ܓ��,J!� �X�۹߳B��tH֞ڏ�R��/������0�;-l-WM�j�!͢��+
�Ԏ��D��Ͻ���@N����N�,�NU�f/=w8�}��P5�x�����fC.WT�u9�KxM.���"���P�U~n�kdS�W]:pw9i��3�|ݚ�,�6��C����i�NH�����c�p��@S�'���>�7�L<+D)��hS���ֺ.�8H�����ҤU�Ǵ��8qu��v ��w��~����=Θ��F6�|��H<eږS^����VD�'e�Kr�?�b�!�PPѠFy��`�]�Q�(�9�F�|��������e(��'��@�ߟ=qw��9R�̟hK"�����iIS:�������X����Jߟ�2��BVj��eu����Rz­e ��f@UT%ۡmK�T�2k�e��%7&���ʩmo��dnf�12vE?%��}_' .Y�;޵�9�upT�ؑ˥6rP��e�R�R�b��c�3�%���+.�m���T?�8��*�h��u2꺶p��;�$��I7����Ä�?j�$��D��;% �
З�� ��7P�-,NA���e���YbN5�]l8�w�\�%�rRo�94��������KJx2v�.���&����Dˢ+�XI�%�<2a��%�ZO��P�޼���]�)w׽�g\�as$��T5	��Sz��}��P�9@���t6�6��Y���T�;��w�e�'E�N������I�/�u�}:I�/�{�zX<U� �u�v��`<�q^�U.W��V+��%�Iδk�}�k./)�Wq�د��K�Ѥp��Dn;��A�D!8x����ң4��`{�e��i�-�J�]$���YEK�2�pͮ�q������rSB��h:˺���ʹ�Ռ��0��� &����7?MK p����Rjy-��I�p����K�������}�v��0�I8'R���x#.�LعWk}4�i���g-8EG�����;���X4X��F���2��� %���A;�갶�0]_���'1I��T��&��)?h0�e�5e�i{��ʧEk�h@���C-HLw�	� �,LJ<�p@��y0R�3P��*��f�~�/�V�M����o�3G��{���L��;D����y�J_.3g)Q'8D�(D�џ\O9��$��[Ώ��T��`YA��dP��N.7���G��'�;���B��<�H��I5'q���,��3JJ�+�RHܴhȽ1,N�IU���?k�AR�i/��Б���0�WV��\���w�O�+�3��`g��ֿ5�O��&�_I�mΡ��)x仝��y���|T�� ��B;�RJ�0N��b~zB�CZ^&d������!��U���|�rdh��8���
Y������,�v��l�N�.�~(�μc��Qe�=���8=��нz�J8֟�l�Z�g�2+�NP0E�^���C�)vdY�U��p[m��9�s�h|��6��!v5Bw�W�I����/�
�����W�|TԬe+���&�ܻ��Y�g����&�)K$��<������� ����Z�S�����@!KP��v�@�Pa:�b>U�H#,��gˑ8������6��=��t**)���b`v���4M,$r��D���*���:��s$��bх-�_��3�p�(�fsAgF�_�A]�`ճ5cq�P��u������ߢ�����{"��Ņ��yB����
E�?ȩ>r��'1+c|?ٰC�Ql�=V��'��M�'1��+W�baA�Ғ)��xy�uN��E�&1M���y�vD͟e9.�9@D2�ЗJ$'�jN{F��_5���?%gڽ$}���z�v&����>���J�a_�]{����_����0ʇ���^���;XC��8d�|�x���V��s�?��K<.��\�22;�G&@ր�Ȭz�iB2��r�� X�t�X��x�R)Go3u*K�źM�>5A�_4t�L��-�Y�����P�-"��B�iڮ�EY��Z�Q���� g��I|T��a/D����t;%cR$�4٫Qi���2M�W���;,�.K���@�<l	����c%Ɩ���C���+ǋ����L=f�Pa8)W��0t�
���C��B�&1��.D�,�wz������s���;�M�-Ți>Kc/�G�n_.uu5�I�1�`;Ͳ��6z��@G���� �k�i��]����e�s�k�V���Aҁ���d�$�Z���96��Z�q��OO�}�W������	�I�Ɩnw@��� � Ru?FIF��I����Q�J$��K՚`@�J���\Ua7�-歠�W��k��0�a�|Q�Vu.��Xag#��A�;��\̿�,
T*�oIw��ȏHn2�}';ɚ��T��3:ȯ�9���Y%�y����k��L)f<R�F�_d���|��[{��\w��Á}a����u��Zsd��-��^��h�x�@��1f��]�b=7R�@���{fA��SF*���N�Ԯ����싵��HE����֮��l	*��L�5d�F��O<�3sbC6���x��j�� ��1���������E�ىQ���*^Q���R���S�ی� ��0���4� E����[�����J��"B���k?�b}��y{06�9�<�d��ce��a��<,+ܷ����&�RBB�=Q*���}L�q
�}�:g!���9�h]�DfjGIF���gb��c��l����X��%*���9�7������,�RƱ��T6���6P���xf:���{�H2��>��74���իj3ktq�~���}5���<�e�?�i�vw�2e�vVa�:$̟Z�&�����@^�0��S���R����Y9��`��Y�4�#����❠�r�%�~���q�W��$�V��>��o3�'LGLֻ�מ�����F
�����v7��tԳ�d��Y��x�9�b:U�Ύh����Ҍ#
ҐN��������h�U��wg�A�%��`dB��y�/���S��pln3���++ݟNQ�"�Efa���a��5��9�4bc����^�B���{gbc��oHK<��f̈́ǖ�!�jU��>�7�(lU��H�:�}���؂i��Y;ŭV��+�%�� ����Q��4��x#i-�<@��/��3e�oSC8 �����,y�w�������ٙ!T<½N��*�I@����c*��܃K�Y��'6]�k����$�<�@���T���pm����L}Ige�ݙ�s�m��h���sS��p�/�V�|<��ᣖ����UhX�jЃ�Ei@�4I�}!��ȥ �U)z�΢����vM"��}�PƸ�m��uP����ǣ}ϼ#����T�3T�����&e鬒�c������t�v5w;����!�;����+��J	ǏG�+���1@p���	Z