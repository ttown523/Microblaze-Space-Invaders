XlxV64EB    2459     b40�3��9�� ���������zДGQ��A�Ѕ�B��A���H0�'۴�5W���=��oϙw�K��!C�:������0���m��
'K�|��K��D���[��Ŧؾ¹�;�.�]���a$72P����MI��
gnaS�|�.�ȠP0g��]��l9�]9x��$:g�ڊtE3�4�+$�0�����9.�r?"�6�?fi/)�m�[�3�;��Ku�vǇ�\����,�fU`P*sF��.ÂL�KD�1�K@�*&� �T_0? ���Hde^~�q�K�4�P��,v��z���VC~s�]D���/g7S@����L���d�i@�gHF��6���yK��6�W�X����g���G��w�+C@�x��}�} ��c���Di���ʊ@{�h�.@�a
S�M98 ��.�Oi�5�t��kΝ����79�L}L�W�o����	ʂhjE˞�d��w�%��׻�6�m�#�ϗ��_����@��;R����9�:2A�5�tF�$�qЪkG����i.����`@�RQpfR�&��F|���������V���x��I��揊��F*��jD)��a���!�YmFF�v.#֥�P|�$�*�a�2��/v��Ӛ�9jZ_��^ˌd���c}E�tҶ�І����Ƀ��Ä�X��zc�
�SEDu��b6��u��QsE/^�Y��
��j����}�\�@���Vƽ��i=��ܤ��ۓ�J|:O�5�I�U؞W,hXwmS�m&�U�sԚ$�Ϗ/};� xcl�
�������H+�l����pT�9MDq�u_
J=����i�K ���6rM�:7F��H�gZ�vL,���A3p���J��w1�h��1w��K��&�����l�q:� Y�⿬��np�\���}XC%5�ٻ,đ����?��sKn�r��4�ӄ����n���p�/RV�ЃЫ�)|���͎V5kH�ˀ���jߕ�E���T��e�9�(���,H���4:Z��b/z��0ql
s���t�~
�\[��QǺ�;��
�
���č7�]/@�z;��4K�ꧻ�:\9�|Z�	�J0,9bgk������D�\�ޫ ��KG��^��]�K"I�b��94���x��%яRL�m �H7�-U3@��qTMM�jó|d��w9����P.�f~��UK� �1k�2���!IaU��H��	+��낯m���b���I��+Bȷz�e|ﯛ�)�YRc����x�'":أ��c�!�����e�/)���mN��iXZU���N�.P��C̗@Ķٞ�p
-m�hVLlB��:��h�k������nK������ �`��ex1	�s5nE@v$�������W���,�^��j���ެؒ���H���uCc��������"=JB=����pѿj2�v���5�ʪ����57G%�D�XV��#.�m�փ�?,�o�_L�$��ڼ��JߥA`7�NJE'"BƗ ����e6����(+�Nz��m�����˨�l;<�욐�����%�gr?�q]^y��B�S�%�Q97�����.�F��/_���WcR�Ux?#hl��#T���Nh24���Xx�%��3j���me�^�bо�9��`�zG��!ʇ�����?�!�q�S�9�3�R.ޭ��D>��`���~|�4bu>�H �C�:�jA^��0A��j���k{I����W����i[�^� ��|r������	�z����o�2H�wЏ�}�]�橴��_����d�Y�>h;7���:�kÄ�"�@�1�r𕭒�����ry����?�j��0>�t��5M�r ^�b��[�yvZ،sG ��S���0c�L����d7]�62��hA��D�՚�{�%�fI��65�N�z�����P������w�i
��,�)�u�UT����R��7����g-�����d���o�Eu�����qGsR��"y	x6��j.�G���@�p����1i|��1mA���6���+Jذ%�U7B������ڲ�S=c� ��ϰ��傮��xfʋ՛r�=�7���!�?7�KrźT�$�y��������띜�sb���w�
�
�h�R_/�� �r��Va,W§��`����U�h�Ƃ����|�۷���0y	 ?�e.7����p,},�'"Т]!�e�ɷi��L��=�*t�m�l�ȉ�h��r�>��%(�9��hF�<�VS�BW�e}�h�z�6�T�]	G��A��WH.�!�>���ݜ|���F�S0��H�;ʾ�:U;�����t�Ö������e6ۖÉ^����hW�z׌��yIS����t{&���t��t�Db��@�� y�W� [ �:=(�f�8Ԅ�<F�M�I��Z<zX<m�=!��Ar��4V���v+���3p||�����T�� �MM��@�"󵜽��s�>bF`��N :"�[�1�����8phê�o �_��3�J�v��Q��[e@�����6�}Ξ����D��>����,AqYm�-�z�O�"-ȋ�,��,!����lV��p,�Zp�{�^���x�&䉴�0 �1�|?�MC�'E�����C�ԇ#Ɨ�4��.�A���c��zk��Y�=x�=J'Ը��44f��Z8��1�"�d���Z*)]��~J�j�Q����4�e�Ĭk��3DP������FLBoy֧3I�$�-n��H6i�BF%�eNS.`:�eN�vvDV����d*i�zhy�l��9:�Ё�^������#�c�y|�'D�~6��M ���f �����