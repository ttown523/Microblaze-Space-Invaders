XlxV64EB    25e3     ab0r���zb6��g�OXjgz���F�mj/V����}ޝ���:P'�!.��0I#�03�cQ�~��dm��A�����|�yTnϞ��r��K%��3��fҩ�!]1L�8? ��Z��q���� տ� ׀1����>�������L ��j�x������a����2
�;��&�pH�����[M��H!w�F>w���7��J�m-Y^ҕ��̙i���A�uSҮ����l�{NA�D�#"��p���F�.���;#,�p\>���� K��])h��:H��l�؞�w��3n��;�h~[@7-:0uSu��\���%J&k�֑ř���uŷ�Z}�-/��ץ��1��I_�M��Nyx�u,��-�_m$�ї�q�zdpxw̻��#���"M���D�B�6����e���G�� �]PtF��ӷ)�����a��78�~�С����Cρ�M:�وD�����1dL�I�¨P^�z3���I�.�eJg%o*pgl�׌Ly���g��₾��L{�k�{!���L�m�&���(��,��ߗ�Ρ�2��f��'e�I�aJ'o��W6��)~���X3f�æ�h��,�A�KmӔG:�x�k�d�W�q�{�ַ� �'��Q
�5ƃ�s"[��帑n�A�[��m*Xv `��b0��(��G�"T|��]���!����L��������K��wE!4�$����oo�uFjڀ@C�*��h�v��-3��)6�Nq��'���])�p��x�!.�,od���p&5ɽa�:,:�����w. #����t��2�0TXR��)��O�V$W���z�4�_�����S�1X�$F�%m{�[d?}�����^Ԫf�:�6)����@Ʃ�"�|�^"��=
+g��ޘm�wǺ`� ���V^�a �+R(�9���_*H��^U�U�FyA��k,B�� e	1Y9���*d����E6�J���a�T���$hK�����~���5�����џ�����bh�_�b��D������y����B4��`}z/�b���ّ�#�=���ߚ����=��/;�������O��oG��r���{6=��S+Z�gm���>R��Wj��4��,R9y�A�{Gy��{����ޗ1:��<ꦁhX�do��w�Z5�2�u�?���W}z1� �y%��J�����ς�%��f�r�_�-X��F��k �[U���|���6�Oر��<8�~(��M�k��}��9U�F��hJ�.J�����{RR|�M�k 
�e�LṂ���g(pN�!iՂ��8b��X� ǀfD�zV}��N������{���	�����ɓ�8(�O�j�]�'5�'���{=��Tx���SmK�I���K^��E�`�?NH/"d����D_���u���񊧡v^���1Z�F�:� ��7d&b�u@I��+�p�lc��w��<c��ó� �꣎�.CԿ���h��z�<��V��б���ɔ:���ˢE���~��$�M�����t��o|�V=kx3'>x��l:��v;FVv�A��M1(��~BY��#M;z'-�V�~ODzع��jn$��_��(�c�A

βS�a�^�(|�0f+#PYF}2�ߚf~2� 
�� �s8��n��d�qy0?9���mQ��vX�J_ӘHE�i/c�㌠9(�&�f\XRL�;�|�>,�v쵓+�����{ш�	NL:��0��U���۟23V-�)<�Ӛ�ԧ�>����W����-酇m���Z��Yh�Y�����م�˩�	\2� ��D��N��4�&B4\N<��Ɇ��'��o�$t΢`���Ig���b�� �U�� ���c��O�|[
�>�,g�UQ<"eY�6���KuӏF(��x�|�7����l0�"͕�yP��Z�����;G@so1����h��4�M�;h#ʡ������Y2���g;D?���W���پ��[��M�e%�ܻ��402����M@�.�'��[����Ac>�"QJ}Pv��98����JqLy֋iH�˩8�gT�+�9�Ll$d`���D#�ȃ剾+2�.Ȑ�>5M�f&�Ù���^�R�l;���vA\�L�42_�@�
J�!�;��_���ҷ����6����a����9ηb(u�EU?9���﷾�X�����<1��{67e�������t�e��/��'q�"��@<G�+���N�A���z� �9�{�#�i���1��Ѓ�}p��X��u:wdr뤹���)@�����-m�@5�)I�Pg1`�B�p���T2�0��l�uq@Z�j�Aؠ�0� ����NK$�����6W���i`k��m~�d�o� ��M�y\�m�����M��[T��Sۯ
?��1�uF��K�p�)�Ƶ�aĸ�b��b��
(�^�3��E�ϱc@d�3خȚ@B$p,��yj�޲WK`7^==Wwq��^�4�K�9W����h�q,h������3�ւ2h���1����\��ͩ�����fa��6Z�����?�_��؂��������fppA8� ��V�:�@<��d?�bqex*�ho�į�4��ߜ}@@ô�R��d��*s�Y�q��L]ϑ��+��0[�/�`&1̇�:�_D�+���>��r) �*Bn�iHy�E��~�Sx|qr�ѕ�� rP�knIcI