XlxV64EB    4cf1    14a0��~�=̹�8-���7���o���[�끒���'��-�Q�����g���	�����T���Fw�ć��|��+F�LQY��7�c� s`IaP�	#:s4>�c�XT�/��Zz%.�V�'"�a;G^H�Кndw��ӛ���s\�#�����q/
$�s����'v�r�>��A�w��@�����ǧ�����A!��P�[<���-+�F=�t���ݟ4�K	�]yX k�ɝ`$/�����l��F�����I���PVa~̹�z�&�* ��͋�M_O�w
��`����>�Ɵ.�k.1Gw�c5�Y-�u`�`ol�Ku]����������33���PP��/�%A!+0���s�3�<o��(b�$��H��{����y��j�	��X�8T��x8��l��5d���Vl��&�����C@����Y�Z���+t� �}�)E�H��(}U�#E-@t�(
ʍ��fU�m��/9�H0�:z�[��]j��q1��g�C�pfKi?�g��V��ObR)�ԟ�����u��oV��Y������?&��֢=Ņ�`	)�}����O��'ߢ����8�/�+�x#��G� ����+������/��X5z
�0�B��{ْ��[&뇦�V+Y�W����N��>�,�j�	޻�3�1�	G䅭���̩۱���K��/=����..AS�^�r�Y�]���\�۵�C$?�Y[BSޯI�@��\
�A�g�K��E��֋��ٻp��7i���5�9k��k�[�:���[_X0�t`�2V����������� �V�����J�V��?�D� F�K����& �v�D�]ր#�u���<^��ҙb����$O
���ӛl���-���@Vn���l `�t���)�s���(LEkì���*�u�c)M$�E�[<�fc���E���p�ID#5Zh���y�?�������g��A@4}&xF�`����(�a����S�f#H@��RC#o}�����\��I�����%5���#�ĕ��k�op�J}3GaS�����o�X�Jj`6,]�N�l��R��;ܸz<0�P�GJD�ש��kC�����C���Ga�H��v��9i�T5v��$(}�CDڜP�na4�q(��W_G9�I�j��S���}]�.����kv(��x�j��d��S�n�r_�l�t?�n'<��/d�+���*�8o8h�(%И��GƑh2�׽T"b��q9O�7 ��M�js����K����_ ��a!�#ms�G��#��V�
�`�����ۤ��q��r�n�-�� ^��z��`���O�N��P\��d��|Q[�e�Vs�?���Hk��P�P�^?�R&�A�ͼ��e�R��O�W�_4v�cZP�N�q��7~v��Kjq�0�Uw+z�)+�������S���\�����GU�C=��N�L�:�t���`�C��a��գ(}1�*�H���D�GJ2��]P��e��Ɏ
�U���.���Z4�ܢ�L(�!��Kyl�S��G�����>X�w:V*zYV�z��*ѝ��(��Z�3-�.z����Y%��C�����ol��.�*��4���"��������������2�hT���ˠ���֦�Z�#̕��y�HE"~�9�}:iO�\�~gt�h�d>�%�S���@��lL��H�w�T+����B���3��L҅<S=c�4U?�mS���.�H�2I�K���8����;0"�2tk�;����.��ʜ��#]�0�v���;�5	�2X���1&ɳ˥Ѷ��*���"�������G�N[}g2|C�J^�\l 		�{���7ޖ��&R���7����������E�2�Ŏd�|zcs"̀`
��4�/�&2�k���"���`��.�����@��d��L�(�!�+�V�
��_�S;��?��w��$�e���W�K�2V�u>�i"I䁈b�����]��)?�
+�U0X \|� _�
K5�VG���`���mu��@�`	��<���7@β�����N��AZ���%�;,��q~��y���H�e��-��4n�K32��VOhS
/�J��ղ���p<�TwyԻT_/�]�Vz�H
��ɛX���
/]:�JŔ�������M�02��ƾ�y@
J9�!^��N�BF�l;��c�u$�8��#7�
���\�	}OF�s�T�_���=��t�(R�b���KUI�������:�8�}IB�<�.;�L%��#��ȾhGZ	ma;"SW�1}�_�%����r���4��=!J�w�6������"$ֆ����q!�y�s��,��	�5�[�"~|�ƅy�_�����<v���(n��.Q��қەkj�,��������`�8��&8_1:�r�.$+�*����z&����H�h�'>�>{��4�Ӭh��r$�])�'��:����g��]:�Ճ
(J;l�fJ�ڜ�W�����T�sa�Z_G2�tߤ~��p�mķ�N��=�ux�P~���[�0v/�/y>�`�Í*���h9�`|�&E 4������̖�9�`��@��6�x��k�xAA�gh���WCZ��C�&�4���@L�g5`9�����Gf"����s�%�i�F�O��G.�����(��; /�� �u5��t�����[*��@��qD�J��ߋn�@��밝���FߴRhc�^�Ao�ކ��������������җ��� ��\����SC�?uX`�;�"^�'�o^��NH�X_)e%���F�+fV>�B��#N,��Y�'/��a$��� W2�h/��*�U�[#'����Y���T��B,qO f��.���'u�|�BL,Z�լ2���9}�����ۆ�	[��e"��$����B-[�UƟŕ��+F�͟fq��ozP��T,��LL���ix5t��1���;�2~1usېd��c{�G+���*B�#���E��5x�;��^�O||9.{�ӝ띏
�o0�5�
;�QonFF�MJ7v�|*�U�i�8��Le5��Y%w�I��<S�r��g��ĭ�1�lpG�^kg�M�2���6�ЈC�RB��⚷�$:�`b˅6�%��5����@2�w�j����B1���<x�.�#�����m�l ����[5��	!n�T�u��0^�]_���(|������7H�y���'_�k��4}*th��0�#)7�w*����gaB'���4!����|�"Q:C�z˲�ea)'�oO	���p���/�]-ݘ�A��N���%�[]�ӑ��( srȿ7��6]P�`M]?|����c&HY�-��û��~�>�u����"��V��	�z���Z^I^�G�ؒ/3�k�w#ܪ����q�N�E�TW�����Bz2�2#����?y^�,ph����d�o^+(�r�aW;�lɛ!O�ϵM9.RsX#J>f��!�҃y��<��C_;V�'�)4p�jz��93��p&����9��l��<Gቪ;(���rtɟA����l�>���n�G�2��H����Ȇ�O|���Kp�1�Ls�9����얎�J)�!f\b�d���K%H��V!d�o�]�Ƈ��ܛ}�K����e�z����´T����ϧ�L���@��B{��YגXj� �]�ZCAVFm{�*��C?�غ����,W���EeE��{\��*L�V���'t��dC��5�ӵ#g�{��8� �R�kw.�EZt�H��g�f��>�t���9�Q�6W�qn�f��ldst �EBQjA��u�S���B����]ê@�mð��۾��>�#�͐+�M��TE��e���\N�w�h����M�咸_�r�ס�%D���r��
)��"����g��QR��e�P�s�!�Mxq�ɶL��g��J��L�{�pV��+�8���ʐ�X������3?��7nN"L�X�g� nP�Z���L�>���%�P�jV����j[�e/!���l�H��Ͻ��C��2ac�E��l@�?O&�My�e�j5�i*.�f�м�!6t��6�G{��[�Q�% �S��[%s��v, ���q���|L�Ď�V���6@��A��Ϗ$�0傱;����D��q�}M�cJ�V��]��h�`��`
���Y���S)�4�#�Y��;+�R5��4��qs�\�Q*	d�-����U�[t��xwxG,�1-�J��Ѡ�H�-4��Uh�.�fVG���lSi1�m@��\]R4��\f�Y�B5�`=�������iiC�̙�X[%b���}�6X��ަό>�
 ��� �{��P�=�!x�Ard�0�8�۩bp�7J ��f�ܞ⤵��=T:/{���3��l��S8
���Đ����!��UZ�/�i�DY�XGC;o�y,��vDros��0���ll���X����	�m�z��A�=��u�X�}%���=�<at,󃴅����_��`�Lk��2k����QeF�m3��)��\v��U���ũ�KѪ��ے��TN'��g�^?6�����C/>���V(��o��f�&�.�;�LV����$�2���D�[0�J���Y�' }'�oϹ��9��Y��G�/�V�`N�w�.e7y�R��KcK��ײ%�Eɰ�����4�C�J�ǡ���|��+:.�9f����{ �Ee�#�ձ�ގ�-!�	���E�X�.We�eq'�! }�%poǃEsg�U~e�+�V�������
;?�x���ۮ��y�99!E�#��)5�%�3��,���g�v��L�_���p~�a��$#!�ߕn���8�tWz�q���9��c���������s�}:����կ
��)na��J��S �L2Tϳ6�X����=s�够1���-zd�O��ޗ�����3�Rs�Vnl	DX�k���&6��NJs�9]�e�B�/���QJ;�DX'��� #A�8���ٝ��7ut�W�� ��T��Q��@�멼<.𧌑���t1�OuP`!�t$��Bb<��#�r�f\.���xo�Rh�fB|�-	�O���D:���`�CU?:���dA� ����KŌ_óa��;6{.�>ga�N�)d��c��g���[�<���$n/ڼ�\f�����ĥ����g���ǚ-5���,��?�[�.�(���N7