XlxV64EB    2139     ad0��k\1����}q!W7	�J���(��=�C/�B����hf1����"�{�f
=1S/e�t݃N����@��^��T� {ȉ���/l�ߋ�}̤Y�A��qa�63�JtU��wa�>��>>�c�pa�<�\2�'�2k��U�~_���ot�t�rю��4�w>D�G��9��l볁SQQ�����ϳ�y����ů�z�b�d
��?�1��5�(���ù$�x貂������YiA�E��e�@e�N	�]ם�T�-7�!��.��Ye���T?Co>ɤ1��Pn.+��NC��x74��D�.��+^N��2Lh,]���ȕ�\͆ ;�q�+TJ8y��7/�s��C6nAk�ŔSQ���ƏtM�O�i�mcF;���l�b���<~:��l���ۙ�h���U����N���|���X~������y���R0R8�}��"�����
Bxl��~<i1�sdZ�m�U3�ד Og ��*}h�\+4���(=P}jյJd��T���V�}��`sR0p'�Ak�j�2s�*��=�3�S��k;���������96Ēh5[���l B-���w�e�<�~K�ӄ|���GG�~|Vz�?��K[:Ə�+.�V��{�CuMjn�!�j��ݗ^�S�6��g��A�>a�+߂+��{���3�ȨKAVm��"y�V��� z3g�	�Y�P��-E���n���;�������j��*x�����&(YRWϼC��'>�]����R� ܢ����e��� ��a�*�{uA��|H&�W�Yi>%j���˽G����$gc�X���Yk FXZ�g�}Hp}l1{�O��?Bk� �S6*���"����t �쌶��j��D/e.;���g�zc;��_Ttq#%[����l�B�Z��Ϲ܇5O��Na9�����M�F�Z�\>���bR�L��y�i/X'�c��<c���>�0��`�=4��~��������j��r]ie����^�<n�G���x�T�=iB/w0�C��E[v�e퇪�����G����"��'�tdP�TX�u�rW��"��X�ċ:-p���;]��6�$��Ch|�e�ؓW
Jഭ+��rV
��&Y��0�@�V�)V���*mNiE���N�.����59��B9��cC^a6��O��u���Q[�q?�p��l5}v��o���k��झ7���&Y��
w�@�ē�⍼��k��$�Xփ� ���z������!�{���ogeбl?	�Ѯ���&��Ӽ�M��w������0�PD�զ��ۗ�(��66��!>�8izt�mir��R�����cӲ�N'��l�P�B:\R�)!)�ʳK阬6���aj������ԫ(V
5ݩ��F�T��̑�����>i�
�	C��}���^�}H�cp�n�J\��������(`�0�kIҟ2� U*^�ǣ��8�K,�&p+:o��taہ��/�Ն��������ۙF����E��د5
��LR*Si��g�hX�P������8��-�ⵙl�vr$u�+@�v~~~Y�ʿ��@����eg++��WG��XS����iWl�#�9��lgVϋ����Y��?������*�s���E��k���`v�m*Ҧ4M˫��"�R�� �2������:jH�C���)`�74QԀ�4E��󋉤Pʈ+��	^J�ѻ�(0�����S��c<�����6�Hu`�[����q�*f��~�\/nR��Y ˸m�@��_a�mX��tA�Y#9��l߿�g��NE��5�t4�2Y{��m���y`O��:��\u6�jvu��)	{K*��Y��3�fӨ���� 锴�k&E7f;�b�a]�х+4AI�&�%76w��Iʝ�O�%�Au�r`���1��&W��ހ��dG�Q�:Y]H�ԣ]	3{ʹ�(�0�!s����HZi��yɪ%y��	����ɯ<�YB���DY��K�������4�Fⲳ�n�+W�1��Js��W�@��#E�4�:
P��{��-�`��ih�k
��^�{�L8^6�V�䗱a����>YB{��bD�����Dt5��u"��F�S����e����pq�X��dr�n���95�K��e����q��l�=6koȘ2
����\�sZǑq��k���i�a�t�Q8�{����S��V0X`ݔ
�����K���jҰ�jˬw/oi�%�x�V�
�hoϐ�l��z5=(�����$�}�Z��]�y��v�+��0��WV�x�QG蚃QM:����ul����@�|�,#� ]L�����jE;���e��M=�L0�H�U��2���9&dPMh��e��ٝ攳lI�I; �wg�.g�X=K�撁#���:F�>�*AK{I�I�V��.����������y�$�"���4J_�5�r�}��L��{9 �4ݞt�5�%�{{�7�̙�Մ�������{���V���{Ј���<����3�Dj'�&H��y|DG���t��GV�A;z�qZ�n9���1-Q�+���֬���?��J�����"����)\avZ�q��0���M�GE�["���Y,"���>�Ë�sM� �����M@c�O�x�?��~�WƗESتT�lph�T�B���U�,��̢ۛ߱�8�d�җAK�ޖ
��U�@s���c5�z>�d�Dp�#�<x�n