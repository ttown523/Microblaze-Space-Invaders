XlxV64EB    b947    2390���(���(8ZY�Зv����e|��e����2D���Q���J�7��KL"����Q�I}4�n�r��51�}s�� d�(M�׺��w��~S?H/l�E��^����f�`�4�����M@��֔��	�N����)��8�T'��֯����^oD�E�k�C����Z����A� �-�:-`�����,�mAf/=�lŲ�<� ��7��6�QB�f�:bE�]呩�xƷ3��˱����_a����Qh\��rL�Իo-��0ق�2��Q+�1���J�]��xw4{��C���sl�G�]�2�o`���ހ�z0�ֶn��cC��?^Vh��]%�Ţf^���C�Cx���AeOVh�����*��D���jU��_�BKw�H!+����	�]0�"aV7�79Z7�����D�hZ�J�`��"�M��Vy=�A5��yS��"/N��2*k�!n�l)�H��%CG��uZ�	�&0�8��x{*����E]���y/@C�l3j��h����%
�ǲ�A���w]�Z5:�ř1��g��TF�q,�G�[͔h�pu#�v~%UA��x;�8��Ģ<3�TU/[��39�c��"������>������|6h�#qIeY�K�O�p3���RdM�Ef��}���o�E���yM�����
7���6��q�n�[U��E��9���R� U�pnL�I;�޼�(�X�����'S/M�'u~�gZ
�4�!U{�����K���צ�o.�l ����[���e��'�4vH�I9k~�X���~;{ꨐjM��|ޅe��? %�3���\���@[-��al�e�l�xB<�X�4� ��Ch��(��lj�W�'�S�>!�oG��u
Q�y2S�Q�\���r�?dOB��������ƭ���F/v�IQL������t�f#70�������G'���/�ަ������=�M���ג�!�e�}���"	y5�%{+�`	}�ı��l�Ւ�2�q-��@�]���/L�?['45-����[�҂C@;5�2������L}	�"�~-}#�Z+�\a�P#W���W��cI�W�ɰpm�Ki�;7�X/�I�{-��k��W3{R�˔�$#&�[;�S� �/���c�t^�֖+�:cŁV8�y#���K�d�0�>����=_9�#����P����=˧6��T,�����v��0q��_2x"G�>h§��l鳊	4w_�,_�1(��0��ɽ�H(���6���vL�0��h���=�Wò���9S��r�-T�g�����U��_˥���3� )j!w���p>��E�)sO���p�T'��[CT
_2[���at>'����6m�ϔ&$�㜓m��^dѱ=�"��g2]����_�c*�T��OmF��A�N]������ܵ��PbN��C� �v���M��@ � �?%j. pg�~����X���j�X��DĽ�C�@2��������>�+�SM�>Oy�yA�����\rp��!��'�G�n�2�k����.*�2��s��ܰ��Yl��Vn��R�H�~�ZN�Db��X=L�5�~`�p�yd	�8!�V�'3:�_)Brm��P���חRi
UCu�ٙ�C_N���v'C�($˻ڥ�y��΢p: ���9jp�F��Ƹު��9�}��	u�����%FA��%w7@:�4��XW��D��Eg�����,���=́X|[mU����j�E~H�}����2N�;L�̎T���OX��y��~�]��~
�ZlJc�r_����J��#	�.�@�y44�?F?��駑,�;P쁟P�+@R�:��c��BߵtWf?�5�����[�|�d{�iJ�������j��:;�!Ă7��"3�\��)lrv��p\�f]�	qP����:�\>�/D��3���l�%a��3�M�fG�W!Y�R"�LS헆�����^E�=�}�z��1����C��� h�ez�EvX�x��~��Lv������lK1~,ɕ�K������zk��ё��.��]��`/�|����f��ë��Y({��3�٫Iw����}�-_l�Ti���H�T	5Fs�C�L�:mШ���A���e<ܛ(65���,�aR��[�!�.Cf�8�bgH��/S�{��K�N��Sŀ�~��]�wd3���#����2!0�a�͝Y��r�vqu�~�a8�����y��{���P�S�0ot���l�:o��y�8 �t����1�U�"kGL�ƥ��t#S'�^6��slOh)�/���<��r��X���xP�����	���X'�8h��28�V��Ē,���*)tc~lܻX-��q�e���e	:C9Ȗ<��to6����g3EEK^�lM���o�o����b�j�L]����D���T��v}]BR6���>
M�����Mv;#"`}(��gE���d����̟+E��/ˑPO�o�Y��S9�퍋l��Ȯ�dR�
X!+�Z�@�}滍��!�Wצ�7̆�L�j�̰����u�{�\���bT5�>5���H�`��gM��c�M���~�c&1<��k���'9����$Z�#O>�0���o<kןO��~�#p
�:��Skp0�6�Ǳ^��0�LR�mX���Z�F7�����]�7�o[��@��
��b�i����	:�HW7� 0�d�OCfJH=��)3�P������>�,60g�˲6�%3���"�6���<�R�Z�{L�hgvhr��X�WAy.�oww�e"tc��)O�R��Ӓv��w�Ga���x�����W/ [�'��e9����ؙv����C��n��Y�A胹���v�ky��v��naȁS8]wK|E�w}�X���$���F��9��,ׯ�1�Լ��AD��Xav�6Y��>�*���r��5N0x7�s֯D��Oi��� r���V��)����`��8GDY�U^�[Z]� ���杕e�yw��O]�Z[�F.�]\�60�!K1VMGg�\ɂ��Aq���Įn�\a[I����W��Ekз��!�e޼C�ǻ�QzfD�jΛj��?�#��?eq�g6?9 ��|"<�a��� Ǟ��"=۶:褭��$��ڮ���)���#)n���G��,J>��%,t�՞���5bUj��&?�F���+J�z��<a$\C@��v���{g}S�Ҩ��H@�Vh	�0�<T���Qw(<	ը�>=�
�X1���-W��T1R��s?P+��{A7dy�������JϏ�]ږu<Q�Fߒ���v�V�d�>>
 T��8R"��}�W�iO��������
V�-�\��~slˊ�D`�1XC���v��Fh (�@!k�՟D�nW,QV�T(��4ý� �:��-�~�Z,2����*�UDn�x�r���B|e��R�c��%�OS�J�L|`LU�'(�p�j��ǋ<"�c����K��H"eDsɺ�3�,gqv����F��8�м�o۪����9*��ղ�7���o�ݬ��=P�=����A�調�2��ּZs*ik�����M:I���G��*g鶠%;G�o�D�W~?��
�Kܜ�
����gO2��a�D��>D�ВP%�$@��������?1�d�v��q��j�]?��M9�łm~���B%�L� �?�ֶ���y��̧�W��Ҝ\�+�Bs��vs�WY�����w��G�qC4ۉ����٘tn	��|DA�	��� )�z2���?��l ��c� mI_px3���"��_XN���k˲���&l�d�����Q^n�։�S���HuS��j������D���k
WŴ�e�}W�����Q�y����,E�Ξ�>${���B���L1�uӝ�T�K�	��Ö(�Etܦ&:{kKM���j�^���E���iK���Nga#�݁��N[�6�2���t���?�͜����f7CR�Q\�̣��QS�F�9�ݕN��^.vj�~�g9�/�t�p�WO;o�\!ܦ7�7�;����B�D�A��5�7���9,y d������#�?���ن6�7�jl�6E�(���P!��D��Sx iq�A���G'��X@�9"�W_�X����p\	)�#-�M�3`.?�o3��F�D�K�]g�N�M�tW'R-,z�r^�(���f�ND]�f�2�S�[x
9��>)�0K+-D��b�m�f���#b|vN�K-R��-�\=����X���J��)6zll냇�v���	kY��Qe�!�@O/��������l��_��:ʊ�$V���f�[��
ru���Ёx��.�~�k^�/�1
>/Af�Q]�jT�����U �Y��"ֳ�O0+�xD�)9��{�p��D���]2c^�����,h�<���M'�Z�Tق���x���6֎�.K�ij�8��e9�-N�ٹ)�j�v�&�
o��HU�;��w"��nVK�Z���v�q��ˀ�_T!���a#$d��j��	�j����]�\�ٖoSK�ֻ���� �BBG�j]X[fq`���#��!?�}��n�Ĳ~ �`o��å���g=-h"��%�����۰2����(��_�Į��bt���ߘ^k01jm�w�����V��,@�c~�� }}�o��(��!繓KjtȻ�&�m�o�󹽪�hf���zc��e��1�)��j����JpI�?gO�͌�kP�lS����I�2����F�NV�� p~s(��U��w&p���]���P
H`�0;U�\5|pȁO5|���r1��΁a�ƅ�t�3*b�~���LM��g:d�8T��gC{J�{�#`t��'�-�����]�ȉtb�ڝ��FG�^c�Sm+�Yd"�ŗZ����D
꼌�D�Ì\j�j�	�����D�ŃÚ���%ʟ`ne1|�#J�c�r�]s�"1v9�j���I۔����|u��*�CN�a��Û3N)X����=o�}���̭�6�͸$ )a�1v��ҁ8�x�V�:\����QX���<t=�;�c�l�)�#�:J���sow;4Hto�sdQ ��M�~#����r�-��Ct&��� �uB�~�^��$�����0�����$'�a���&��:�_3Ri 6i*P�r��Ij�$�|Y��bm���G�^�O*������3jD����	PR|�w��gP�}_�֫�� ��:*+`b�Y�|G�[��h�������d*4�K@�0����RA��wF�i���xe�i��1Ǟ0d,XT�n����XF���kvUi�0���@K��`K��4�ڴ{�y$�Y'{%:�U����.���r�D�d,رҬ�S��%���Z�\7� �ڀ��D�#�`?e����ObE��t�|���o�����1iN��`ay2���^#����P���)�?�ڹ�"�{(��G-����xjjV-+�)]p�z�w/��S��­K:w0�+ֻ�T�'w��/v�`r��T8���]F��/� 7��"��}���h��m��>O��l�:7D����g��Gv(>͟��qy
_��[��=�KM��wÛ8���i#2;���b�,�^��<��+b����𷏀v�� �˻���Y>r���Ԏ�9�+~(�խԳU�W#{S�t���L
�ak��`�;�Mo�� �,������Hy����������^�[d$�	*��#ӈ_N7ŸN;�PF����^�>\�y
eh�r<�U���o�GWdY���Z)��B9�`��`xa��m�j��&�t�`���1�y�D��JC띶O�N\zW{�EDqgvw�s ��t�&�`!u#����0�0g����kW�� ���K�_��ICv|bnj=���G�uH0G
��y8�q�L��b�{�*�ƶ�h��ٹ�d�"�ꮪ>�(��m��@�F�����+�ݷ�N�����@*��<��!(i�x�b �^��d���Æ��+�o�X�����5�A��Ekr�ji1vq!���W�;��A�ef��˫�Ѽ��J ��e Ed�S��"=T�SOS��].��.�V�&�^݊m��f>������ƾ|��۪�'�o�,.�S3jk|8�&����9&7��_��u�4���3C��F�s�_��5J����F���;,�����[Y5=qv�h\;�X��,��Y_�lOKV�rLz��CY�;d���� �F�/�WEq���v<��M<���6.� Ǆ�U���+����x�$ۓ�n@�։���HcI��1���^~C��'�¯)���\J�ms:���e�W+���r�w��	�*�KL-���C�̟����XEǰgc���o�΋�u��em�r煦V98���-�6�
�������ri%x�<���R'��$*.��%<�ohǚ����̔>er�O֤�:��	2���X��Y��)������"#d��}��1����ĉM�-'=���s�Mtć��3�q��,"��P��}2������)i�!l�@��)�2x���gg�I���_��b�)&��t���$�ŀ��w#0��M�OH���}���Y+�j�9�������Wc�a������'A�O�ok�J�̰TZ����

hV6����aT^� �� Ѝ�(�+o$3����Nkd�\D]A
J���c"q/9���tr/-DJ�(���v�[1��&�ڸ
߯2
�W�g�2��Nzv���%~����&B�m'���ؚ<T�	��<4����-j}����"�8��J� 6�1�p�U��};�W���Zw�o��bH?5􉦜��#��.QLxޜ�ü�U��'7�y\s�^t��PٵUlb��}�1&ČLc�y���]d��5,��ɏ�r�#B�Y��⹏�O ���SK��f������� 8�� �6��2U�0�ʵ���̄�	:G��Ű�?_�m=�{��rDVUQ�H��3���4O�9k�ߨًVy>�& E���c5|G����\���s��Re�Ch�ӻ����wc2��w�su�:@q߮j�G�V���G*�+�M"v���_��i���~M��>���˧2#� ����)۰aC�����%���}���-���	?���$J�q$�&�恇�6�N��o��U�ۂˢ���w��S����D�xj�dG�«�>GW�~ݎ�5�ziJ ӈ���+Lٸ�'ˆ?�J�.+�"��g4Z+�/�&T�%A�͹�L����4�0[aA|�U`c�@���$;y6+�U�Ä���MW�;@>�+)�g����6|I��a�E���:WM���s���, X��W;]9w �]�p�0a���=����@��I�����}���Ԙ5a캢�[D��,�HqB��Fy[.��l�K}4eI5�tM��|�{��G�8]Iv�t$�S-�}�?Һm�vG�T�ᆗ��Z_�舧�F;H�hlA2��E]c{tnP�;�O�3������j��|�w��=��V���vqSD������@���5GE�lF�Ql}�D�v"��۔����Sm��6؊[�׉�fg�4���\#a>pP�ͩ;0Iy�����h���.D��1�*��@�_VeR`؍�qk�xg�;=�\�U�h����E�k!�MX�&s�Wx��0���\��]��O*��7��~��MN������/��n<;2qd��/^Wi����pl�4�wR�㹫[��p�i���s���TE^ģp���\��Ԗ���d=�b\*��e�1�6��^�d�Nԍ~��3燦uؠ��݊\�?�$����[SRD�����P+�T�x��@Nh�1�,�8Y̕�0d==K��^K�˷O�i�n�j�%�oZ
m��^�Jcj�3�t*�����R:�Y��@֒����u�;A��Z��?�+���f	`����5X+C�S����5��>:��>���T/��-ЩA�"GG�^��,�m��:g� ���& ����
��f���86Z�-��c�\�iz.C~g�ZA`ѭN�E>�b5Q�h���D�i�K �W?�O,+/}5�.WsU�����L+c�r1���ZQ?z��k�?�j)�ު�Sg,Ɂ?`��.��:@ᥐ�ɐ��&��-6�@�9C/�%'�y��<�/��tL�����F��9���aj�C�a������ϫ4c�fD2U�Om�0I�D?�|c�v��}q��v�W�
��=��\ š_��r�f���J�4���O�n��$l����#�;N
����H(���6E�ЌJh��ַ���N�W���L����D{Rjx���K_c/�[W8�щ� ���q��-N���R��0��M����椣t��w�}s/��{M�E����U19����*衍�o_�j�0�h��Z�V��MJ$�ƃ�.���X���s�=H%=��g� t�X9��i���\�B�ha��[]�����楧Wv�A�;d�I#T X�����>���l��u$�~(�D7�f�ܮ`�
�����:ϫ��@��ג%�>ۓ�5�}(nWI@��LōKV��C�7CN�����0b�7�5`�
(Ъ���}oK����t{F����;�1�o�|�{�'�
#�����"�x?X$��3�����OŽ�R�p�#yO}�i�$��P��DG��U�u����a�u�3ـiX^-��WֳMo�����+�x��o#�ER�n��[O'e����.��u�K��?��+�Bg�ҫ�>$*���X�R���y|�Yu���š���Xȁ2�D���w�d�ټ
%)�`s�+�뀴��g�r%B�)���\�9�A�k��K���}r�	�膸��)OW�e���*���i ,�Q���`�qJ�S�#Ӿt��L܈�舡D�5��X�7/�JS���: ���`'�	��S��I��%�>�W�Ǩ�t���=��g