XlxV64EB    162c     6a0�^Bc��A2�"Q��&s��bfk)F+�Ƴ�z�FSA0P���湱dY�[�)�{�+W��}��
�����6��6~B߰c*�4��|>fxjs�'��{�D�t�����A�ϸ�y�%A�x��LӶ�_��[�F���V��I�og��|�u�İ O���m���u[@	&}4�J�ʭ#Fjr��[��a}_��G�Ȳ�c9Lu��N��'Y�]�����k�ʟ������ז��~`� ��`��_���@Ѳ*m��xnv��M=JyJ:uFM���w��Վ��vs��$u|fz"�����9��Ҳ��C�[d���V[ڤA�޼�1a���@�x8��su� ��qUF|>6��Z>/K�K�'�%\�_Z�'�}O��C�rlG�o�V��(+D�	`�[�v%�)X7L�L�����B[�oi��7^e�r��P�g�9� L����?7�2@^�>�h�v4a�"�Y�Uʴ� h4�����v۝�MZ��\.�U�F�i����-���я��@�Ȗ{S��Q.�+Lx+��K��Z^7��2�>��rZ��Y��eʄ �<r��#��Ħ�j��+l��&��<��7���v4� ݕ��Ƀ\�f|���ſ
�b�w����aa�m�����
~]r����{ۊ�Q�ִbm��زN�G��h��@b�]zwo;_�\L,:x�C|r�W�-��=a������Ұ��j��N�:%]k����z�j�E�W��z�<�H.j��e-5�<����p��{�jH��dc��}]F��G-#=��p�ȕ�����&P���Ȼ�E��8��s���M�O��u���(l�9����ؚ���T��Ԅ&�d�]*R��|=�z}��S��iC���~ԑ-݋9�*�U'�������^�K�%��$r��%\�"�c:Ɠ�F�$��� z�s�!F_�^tS�� ���o����H�hݭ���EB/	�0C�e�_a��Dh�J��
tZ�X@��	)����"��d{��������g�����<��%�F�����:]�P8��24$�P��rSż�s���Efv�~h��r�Y�4��O�2��� s}_c��p3$}p����lp����E�6S�{�
�A�V]Ҟ�CG��(��v�k�.�B�rMc%��p����ԓ��;-Ʋ�7]�];S,eޡ����f[�@��C[wj��\�����>��f��7�+ӂ���|�#�>&�w ,L����tO�dk�u��lq�:����$v�]G�:�/r�Q����\!���D�i,����ɯ�<}�����XSӕޢ�Q�z��a����hP}q+��6����l@M$%	,W��^-TJ�En0@���b�r��&>�c˄��)���)x<]�n�x�ȃ{)�bb׋�iE�v��	����wD=���*R�w�$U�����.����\޽7}����(x�gB��9��u�9ͳ��k��3�`�DA�%'�ջ�!��/F�q@�ETw*JI���7��9$�z=�Ͱh.��%D_��||�E��n
� �uk��]�PA�5
��h�c��|�櫪��Suo�,��ٮ�QԽO=62+����d:�N��I��95-�5�2���u�(x{��y�l��lWX�D��f��t!��W��mo�ks��&�l����Ә���lD>��B�
�7�=i���