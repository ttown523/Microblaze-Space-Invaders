XlxV64EB    187b     8e0�p����<|㓶q�P��J�Y�h
qCg��.����9ڇڶL�Ѱy�݃�z�l�Hg*?���.;[�"X��#��D�S�95*+�`"-=�xǷ��:W���~��Eʅ\;�A��H��/=��7:;��i�S򁯷i�y�i}�|�\̒����O�>y���9|�Ut��`^I2�H��r*��h�o����@�@y).���aW��2Q�' \*�|\����mif%�������LY��Pv45`*�*"��h38���F�b׺;H�|'A�=�1�-:�8R�Z������ҔP#c$���v���lu���JsV0oѓ�΄���L�8HN�����]��1���Ԑ�u-��h�	i�sp�HnI;H�-�_Vu��8���6b�l�v|�V�(ε6a��a�ag����i���`��Qa�R����kԒ�p�o&o�xԥ\����o9��^�#�.Y�Dk�ݪ��P��˷Aq�J���L&&!�}�=��"�C8F ���[{�K�,�JQ�Df39�ف���Ը>Ư$���*��gg��S�+d��媉�p$��;�����H�)�P�y�?�7+�SI��nd���9�X+�R{��/R-X�C�x�+��� /Z���lݪ꺊L�}/���ʄ�Sr�aSr�1�����{r�e"����K�]��]ѣ3��ĘG�
X|	
�{(�� �?��C \,��Lk]4o�N��^-
ԣ9W�ԓ����FV�y�Y����V&E�Ǩ�c��)�6"�e#��c:٣�@\^x�۠��܇���ָüW�}%�ͨ�F��(���� ��G�I�:[2��qtm��s���Ev��T8�/����z��r����Gy����)/��C�� GvJ
���H���bj]&�T<��j�����˭x�#���Ϫm�7/!0!?�:�M�� �3H�G��&�&m�|5�m���}S�
�{�3'>o���
�*�����j��aN���p��W\�W�s��	YH��f9�i���2%�z�to�qv<�z���u>��yp�����y_yP��J�֖Y@��tf�~���&�`{����d/^�4)�A�r1�)�Rs�<õa�)#������O�LV�tho�TM�,�켰iu�}d,�����)��x�P5.�rB�A>�ײw�%/_�>�����?!y����'"c�?h����(��`ǡ�����W/O���rie�q(�0>�ꕭ$*�Na_�xJ�D�ƣn-�ѧ��\�,�o�9A��ə��C��d�B���a ���FŎ�)�*}�ր�	LyJe��V\�G���(�,������4#�BJ�.��@�Hİͤc���L�o�_ύ
V�D�Xt�v�L��%��g�Q١\}���n� s���o��T�������D��춋�r|+�$���#(���MT�F�XAf5�v�L����3�6u���Gy9�}/�E�@�����e�xd@���E��F��6*�>`�7b���'psf:��US��q�� @9�����Ιl�ړ������k���{�P���\
�7kq�����\��U��^H��$JQ��ufhc$�m�/�`��/\�~s�����ZM�f�"�튛 q���uHt�B6�����w�?�]���<��4^���4�^�?6(`��E ���2o#��R���K	`�G��I5!u;��
�⹔���jW��~1_���3E]r���Hkc x���o��T�^�h��]4��fdr.xL5�za[U��p�ø��Άv�j�u�˽�Zz4�N�Μ�=8o�{e|�qg�����u$/P�=$!�����?�-����۹����cNd���+)�$�vQ��e3V.?}lZd��WILj6@mj��H���o��ܻC.�삁���4�������I��65���ZZ:~� 4oHKo{�\b���R�
O�(3�B9yU�&���Y2I�p���ⴰ��>��+퇘�����/��*�#\�J��R��ӫ~����=���b�2�I*�k��~ow�(��8�r� ~�'vހ�aIr�2�,2+�����]��F�&K>��	��Zx�듘8q���Acn��t��B���o��#*&q�jq��<��:�0��|�aTIγ2���p�7��8�V�!�MXtOx���@5�i]~�m�gK�_���됌��Hf����?p��4����Or8x��2�l~U�W�ѫ }������y�hi�Tc�,�֗�