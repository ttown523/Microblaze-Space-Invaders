XlxV64EB    fa00    3010���-���L���'":���L�� ���XQ���gRszG��y�[F.�ި�q�>œ��|O@���:��_iV���o���u��P�-.:ޞ-w��,�J;���m%e�1�`�i��=��g��o��g�?��]xI�1r#|�@|�\����	���0V��v�vψ�>R0�x�J��ڢ�*FCiIѭ��-�Tя��)�*Mv�2.�ec�*����=۳��*a��mʫXW�,�5����=����$,�2�� 8?��fvO�˻x��x^/�?�qSO*[LH���5~�RUqSY\Ap2�0������x�:���>?@R@�cyopߩ;��!]�!?�w�њP�j���&�����$�-���T_���"��G�~6��Vb[���:� �� �Wr����J�G�����O�����K܋ng
ܦl�`0��❊P��8�ǧ?��� d����l#���4��k6�iUyE�q��ԣ��b��Wo@��I���N.z�`�ۚ��$6$��nJ��T �z�v��e�t��χ��*{	�@�?�������c���u�j��$Ȱ(��Z<\ٴ�;�j�r�Df��h��ԤG�Z��$�&��Az��6�X��W��aNB�q��In�-b3�h���Ι[͑�wxFE�~FG7��R�y"��\�(1�Z�Հ�[�96�%�3�t����f?C�ߛ��M�v�1A��ȹئXc�	N/6w�9�N�!�r9�Z�7�M�ɾ�z�®z��$�1lh�rmG8	�0��'���p}�L8ue���+��hˋ��\X��$J����;���Oլ�a��4�'
�Of69R��؊o�)��CU���$dFG�1��Ѓ��y�">�z*F��\������d��Ka�G��YsaT�Rw�&;��"g#,��5�42{.FVߜu��ꆻ{�-�|#u���y����9��cwq�?V���i)����˳��^,�l�"����n[v}�Ei����?J��1��?���3Y�^�j	u��/���=y���k)�Hkԟb̰��
uG���p&��6%d�s
b�_�	�{#��T,r�0�;?��nY݈28u��4�I�<���������g%��s����~29����nľ۔/����,}2�":-�K$��
>���A�	�GVi'!�ӝ��e'��2�{~��?�m�$�jtDC��(�fc��D��ARQ�O�ׯ��I5+	U���k����BP��	ֻw��J���}c"�&��Tq�H�D�^���m��ۋ���T�J93�	� c��}�f.�>K�P�����HC�/�'_�'eG��5�R�(�ק��8�m�>Z�a�uo�,�΂��3acb�Dw�+��O~]�!� ςZ��&�x�Pa�
m����G�ϴa\�m�4�e=�r�L��q����q\����B s�������Cx�rVn����b.�r�x���C�/oM��z��D/��5����bk�u��0��%YJ�?r���>)|��/�f���@eQP��:z��L�lDҗ��a����=�
�Fw*@�b��ۣ��L��&�Ֆ~��"igF��sw��d	�ߐr�<���X�/Zƺ  >D��������U!el�1���\yA�_�u.�%� �B�
�����ĩ"�i����n���Ҵ�d�&`d�Nx�EI����98�ӫ�vZkΡ2���i7	䄸�Bv�ʇx�n�w���2it�7k�e�[,��;6~��
�4����*��c#RN�;*�fK�-�;�$��9󇛝��v��gG�Ga�Ik<��ŁiZ���$�igd���@���iɸX���`-q����T�f��mƁ�����lR��ce���SḺ�THc��K��G��.C��!Wl���+�"%8p��-m�à��Sz(X낰�2�P��,|=PrƲ?g�1!�@+Ov�۸����Rm���f���S�O������PO�i��180XpA�ܥ�y]u�^�e�}7?�]Z�	�[��-�\J��	Ti���kVb�uj���4��<))~��̻]i3��~�C=�7�l� ԑل�.^.�<Ue��7���K��/�����������o2V�A�Y�����-bG�ϼ��.Ԧ���Âj�G(3�P��֨E�`r{s�c˯2II��Y}���a��K�2�1�$TX@�m�+�<ogY}�ɇ~���@���Y@A���7��n�uY�߁x�~[S��H�EoNz��_�Dݶ��U>���Wٹ��N�
�{_��yj��8�]��)Z� ��C��k�yմ �*�R�V��d�����(��Ҕуk����A1ȩ��-�w�@@)����h�$֞%��_WTq�h`���8_�l/��@w5ݣ��y��A�g˨ݘ�JF��T	�f��ڲ����ND���� ��x{��q�f��]Y�$�B7����Di:�_i=ֽ^78~ʼ�
�4<�<f7��nvXpT�.�\h3'�@�Ί��!�J@1��hH��l;����i��+'�ߞ:�4w� ��[ix�rؓ5�ٜ?>r<�k'���Y�\[�L珞��������`��:���V3&��ªOay�!��Hhq�<����>G�#�ciG�S۝���G��8׭T����8���}JO�@)��� ̉3�^dk:H>+�S9�S�k�umՊ��ϬMߐ3(,J<Tv�c�u?G��=�}��t=��u��7;�2��P,�t��L��p$�e�ՙ���Ⱦ��|#+˿p�?��8+�j���Z��U�O{&>��"���T@���g���=-:r|m_ٔG�Q&N��?���T�&�9�(W�8������w�����_��u�Qz���	���>6XoY�l���	ϐ�k2��T
q��/2������l��/���0��6;��D��쁦|9G��ȉ���X���@e��.�~Z��J>�����1�솄���F�7{�q�@)�wI�f*@�Z�7��V���Ǉ��y�����YX���Й��I��#_�({�e��c��� �z�'_W��3
�#����Ski�-�����
KԬr����զ����:�8��0ց(�����MS�>O�3�6��Թ#P`��GO���hx�:i3�g���Q����B��Q��K�h�f����K�́�_
���C|�w��9����3��ޱ�1�K�+��eh���I�����D�>��b�u��i(����-���au�ڬ*��@+���!�F�죙Sh�c�������&m��p!�#چ��r$����ϩ�]GL�({��U5��������B��ٸ���՞���N��;��"t�n�޾��;��9-"�#F<��d�M���ZU�+���*�Y�`���Q!�"3rY��x^���ZOU��ϲ�l]=_�tD8�����g�dݟ݅Ǌ�s�g�)�C�I�E+�	"�3|}����7�pm`�xK	7)��D�M��ϻ[d��Q$�&�$��o�PiF�`6z&������5�HE���	Q$�����g�%悛
R�.�7FZRj�(U�����:���(��?]��_�E�G̏
�`���_`��᜕��ф�Y�P&��������D�ETpJ �dc���/9�0#�p(���iK,���7��,�`�Xg-#q����Ё��QB�5m�l
��xB��c��w@fB�\=�5����{�5)��@���wl;���AY�H��IjE��t9�0ދ���vDr��طp�A�B�p܏}�
^OU��r�A;ST����Avv��R%nP��M�6�F�|�Ӥ%U�z�AwoX鶖Q�`O����J\Oe"�8��6C�wJ�������Ջ#�����?~Acm�U�kF�L�������r�pcEu�"�/WpY 6S�Ipg���1��wT|��T�B��Sδ�)�Ŭ ��MN���Jr�
��[gg��'�hEҢ3G�G�w�
��l��e��Q?���P��w��eAس�r�������Q ����@�UZ�]���5�GCx��/� ��=>x�$�<�=����*}���6#�cR���<���g�8�r�izE��;�}��5z8Ox��&�9�'�JU)��F�m����&����y��������,+�����@�$" �ߺi}����W�C�^�MB?�ʧ��NX��$�C�\T������4K����n���/:c�ug{:�CoO��������D9G.R���t�I}���C��jdڛ�CrI'�N����D�Y[����Y�*�&���D�a�aB��$�|��XV�RdPQZ��X'����$�.'�%�IE^$p���^�1�<7�����NA��Di�n��x59lHGG��,
Ę���C���rւ����Ȋb�����v�]�؇�l����L�-���S%��U��&�I3�'7�'���n7L�;s�(u�}"�բwy䗽��17��i(מ[�A��}a���� ;th݂���.) � �)n����
������d�C*~���qM�TN�B�<��?��1f��M�0�Ӂ�^��H]���R&�qo��Wi~_��;�A�RžwA�=�����&-��ЁL	
����xj���k�~�{��c���k�P�Xy�wL0e�I���3�~4�������O�:���EZGN�˥�8,f@���8��u�w���a#��'nX�q`�f�ժ��M�M*E�kხW<�%1�fcY$�
 T�E�u��I���N��F��~��Aº��)=M	�e�G�����:�$��_'H�*o�lI�X]&�6{����9���"�˦'���T�� �9V*>��e&���ʧx�`��8dب\�����4Ê�d�!�����)�E�ae���!)���g�������d��"2%�L�e���G�|P��s��4��>����Om)��/i)�� �I�\Yk���P�s�~c�������d�9��oU	��I�b��Nuo��8�����	p������"�ǰ�E��9�7%|�F�d׍jS�Bv/��ܪ7�Q|��^�]��%g)oq�f�������N�n#lr�U��s�;���9/�q��w�C��域^2h��G�n��P�n��lP
aiգ�o���`�|t�[D7�����\[�0�gP�r�^_���a/E�?7���9���&K*�}��AL�SFn��c������*��עNҿ���H)o�����^�Oe"��[��>�����~R�E�s�ۉ�9b�	������.�;U|^4�K��Q7�>���(}=�_�J)���<����X�ո6X�S\�{HN���GV�@�{ns)�S�K@�we� �I�X�@A����v��a�_��W����_7%���+56ш8?¤ޥ�\H+c�|��pW�TRV4l�(ك��?��k���٥1S�5��n[y��њ.� �EE���7�b0�)�Tv�C^�Y�uB�%�R��ٙ�Hg���ëϪ��ݒ��E!S��uI{.��ǳ�u� �q�3-��v�>�l��_� � ������<+�����I�Ey|x+o]HX֜J�[��%�?��渢���+�����V�.�:��W�=ߛ��B��+��ap^��܂b�R��V��������n��x�o�ߓ��✕F�+$�e�6߼� K�1���6<m�{�%vh�����gh�xF��bpD�c�gr�a�w:��n���h��%<���8*���C.�
�#u7Ɖce�>zm��m�'~��$s�x➙6f�I�Q1�=Ā���}�7��Y�Dc�@|;G�7
��������'��x[���Z��V�z��|�z�{����J7RRj}@�!���,4N�̀6	d�"��[���G�4^���GٺR-��-ͬ��U���F���*CS��6�.�^�
?e�uH���fÄ?9���w\�K�]j��x��m��z��u������R��)#���U�,,��I�=���xހ��ܮD�z�I���ycl�#wg+�e!��&��fs�f~��W��J�*���7Qp-gT�%$��۩>���Ut^�}w4Zz��Vw���gD�_�ʐS"�ٔ�f?n���M�VKj�|�O��4K&�� 
ϒ�P�f����d���3O�������kq��۝�h����&��g}�Ҫ�	y��3�y�x��ܴF��1i�F��ˆ��3��T	:z�R�[��iS"�M�����9��Ĩ�
�|ʜF�]�6��|ń���������̳��*���[�:"�J�{���Q�ET,�.5s�j�?�^t�3C�J�]�뤇�2�e�ԆR���#��K>��0?R�1��X,���YI���+DT�Cl�&)��LXs�
��#�)�@9���IF��s������O`�G^���h�7�o�&��,�O}^�dI3��G����pHڊ�+�<	�+�N����C�JP�|\!ؕ�[QP5h��T�P��Z67�H����O��th#��u%϶�X⳾�L���:�#����C��%0n ��X�4T��ąs�.�o�a!�"#����8G[5O|���:�H��6��0x�(��vV]�:;�VL�`{$3��$�%0�{����%�wG��fu��Z��b֒�$�WN}�z	8�ھ�[�ߔ<G�Tf��#ߡ4�j�#X=I=�n\%P�(�G��X�l:R�H�4��ľr����D����m��Ȋ`O�g�5��<���;~U蠲f�6x��~h�Yv���Z@��8�g9%�õ�H���Y���l��b��i�+�ӫ�օIh�����b�Ĕ��G�����u���k��*�1%�ƺl�1�JJq�5�h5v{i��KI���i���8�bl��t'�_R�X6�NC`NV�'�ؐ���V���7�n��^(�����kh�@�R.��z ��9�vV��;����R\�sq��2AkO�d��4Է\�^�e�g׎�7���==ƨ��]K���Q|Vn��4��tD}��g���*d�l�@&�^'&�i�9��8l\�O6��)J�����Aؠ�.���t���`�N���bk��Li�9�C� *c[b`F#��z��{_68@)v(־C���JO�"�o7�8u�+o���S
�/^����HbJ��>C�־1Ǉ�'��$��j{�[QiQz��:�Kj�>,��e�95�4��%�P�⡾�������5E/gÂK�;Vx�i�ݜ����g7�l���"m�����[a��E��ͧ�K��;�}e�~X` m�<*�t/���"O�zq'��B���|��M��l�<�K���ۍ���D-��g�#%"����4a��:�̜%0�g��xvE#~��3�sWP9��U7B6E.�<RJ���KÙ.�S�v�Q�(B�=�����F��ڏrP(&��q��{
�Җ���K�H��+P`Gs�=��f/��"i�����)G-�&�~����
,��M[��L�9�kt�Y3&������t:Z�Se�T���[�B�&�mG�p�:�D�0�\/�E>�(��!� *s��7�V��Y� ������u����:���ה%�������Ù���/3yZ��\nv���[�=,�������Uۘ�7Qd�Fuh0;L�UQ�����q�[s���������)�,yXk+��L�����ޘ�G�q��؜>��a�����,���s�Μ�_K=����10��H�8s�oP��������;`չ�",p�Y�ߔ��+i{�U}$�����\J*顮�opЮ�m8�h��n�03�^g�ߜݍҋv��D��w�{��p�q�z��/�)��]&���+ ��G���Y��]�'�<�SB�@�hpS�si`y>�#h	tF���q/N�>*��)i�G�TZ�R� ��	�%(m��.�D$X��p��d�^�08�12�y�Tl�du�X�C�ut6K����_?�E���\�����Ø�ǎ)TX��jF4���j�Qs2���<���!�)��ėɣ �;c4�T���� 4��Ղ��Yf����ZE�f�$�� �t��Ze���-�q�)䯀���t|$�L��K���o�Bs�%��(��I[CcAx�%�vq�!�E�EK���yE8\uj���䗗�/#�C=�+��p6��mc%���NJ)-Q�_cJ�#�j�^t�BE;[�TUĀ��K*Z-f��E�=�:�+7���ī�w���7Ŕ�S�M��l0��DH���Ե0U��xF\�1c)|92�ڃ�JK6�0C@&?�8��^"r�q?��
����i����ۿ�M-��Sy�R�a��蚥�爛0�9L��)ۤc���t�V�ל��*&�+ފ+������v�=�Jށ{���<:������������F^��Sw:'p��S� @OƐ����w[�Ҩ���R�~#1�n5�L���0@E~�;��먦�X����uW�K6��C����nG ]�ګ7Hz|V@�?MF��(,2���E����ۡ^������Mvv<d�# b���7o��a��� ��rr�1n��;����B�_Pc$�����Ľ�g�$j�8�y�ٕjINn��a���|�ٛ�p�X�����&�}:�XI7����{�Ғ���	~����@аi�x��1����B���S=�]�+n�qR1랃B�5�_��hI��K�O"7��t����ϙ,��'���m��X��F9�p&ź�8�H��غ	��R�v'tQ�%����|�Z~(�JC�H
0C4��@�*
P�U��6`J������O%6�����WiP��<�"�<�[:���
h�S�7 q�$YF�ىٸ[����7�C����
�Z"�g�56u�>�3��ޗã^�;��ZvN]L&�����k�#~����؎R!���D��a�6��>C��Ufc�45\|��ψ���&�l�ʥh�L �ۓ,��Z@�N�W��{V��F4�ݛ/���Zu0�Ib&3�6 jDU��N_ਃ�U�8�	kf>\��`Q�,Mj�%��Fe78�	5z$���<G}1T�	׭`c��%��S"��n�Z����Ϸ��k&��J�
C�e��7�q&�TbD#.<K�ٕg.rIU��W\�������ٝ>����aÆp׶iq
l��IA�;����ңzY�%�>�94xf��R����զ�n�~z똆gY��������AC�8ƮC �.b�b��*:1��(��a�_��e�7��GְR�e��S����� c�5�ƤJ�)��	/G���ʎn��z�v����ls�d+�hZ�'��5"�ѹQk7��f9�2��o���h:89a�drX�ʆ��IMfWox*��AYɾ���u4ǚ�\�`��
|sk��'Z5c���aJ�m��l��:<�ą��e��vT�9�e��~�Z�h��j���Ӌ��4�F�o0z ��(����=)��ut�k�$VZ�fz�o
��9��3�����>_�>G�� CV咆ғ�2L��h��A���㧻f��L�T��6��Lt#��^���?���YvV��q 8C�$j��}��7Y��Z�*��a�9���ڰ2>
W/=8P�Q+���)�9b%0V�Ś�b�G�@`�"���Y�jY�a�2J_ܸ��7I|�����B��έBӷ�?z�b7�v��n�Z����s\&�B�y����2����5!%��{Y�4]x�������mБ��Z+�'�Y��!�~��Y��PQ�hEy{�Ԑ�������M
�1,~?.��7��'�NR�YX��?Sq��'�̋�lw4�l�~�w��$bӑ��T�j:d��#�ݩ�WH��J���V��i�^�4���c�g#?��Ѻ�^���ﳄ�E/wL����m|q�źǃ�hJ�@"��w+�O��j����98q<V�ձ4u������6�r�v���lM���
�?����Jºy�-�,����hI�fSIt��?Z���ʏ�3�������@��E.s��p�N�O!*5��̔���슔�f��3�lw��y
;��4f�Y���K�D�!��'���* �'1<�>�Q*�V���C����W�k�H &D�c�ڲ��z
�rZ6�z� ^�ם�(� �I�cd/�������h�$@����Y��~B+bdZ��4؏���!rP4֠�ZoF&y35EJ��w�ļ&B�����\�Z{�ˀf'f<�� M�6�,�6z%���������3��C���ه,M���|��̵�>3�^MUx��0lS��oP|G���w�mD��D�����xnp�
���}��ڬՀ�E�Wٺ����Bp����%6��Cam( xϐ��2����$����}{���#��QM,D��g"��ژ.�ޑۨ1�Y�t~ ��=d��m�Ԩ�ף�O������Lګ�	��b�pn.��3��Q
�L�k%�J���#˛wv����Q�oU3Te0h���H&�Z����~�d�Z[����:�"�~Q��A��k�4a�e��1�0�6�[�Rle�DH�<��!μ8l(̬/��	t��g�؈�]�O�'ak��cfC"_~	����U�ix���W�]�s�E/a}��_�)H_�$�J�������޾��d���n�q4���cb�01GHPP���O+X���G�[���ߓ^�<�x��I1�z��bW��8ͪM$�c_�P��i�_���(�E�0z�M�7�y�݊��qm�b�HHձɺ���E`�Pgr:�h(�Fю�U�+Tg鳞H�OP����1��,�jh,�����;�{�tZ��ў� qsֳ`^�n���B�RV���51���A�kc���D	S��k�V&���!=���|Q����
���N��]wԏ���7� H�o�C�_(ʰ �g���ːnB�,,m�6�|�˨�x`�/s�����v�����+F�NNi��]ÓI�!?��Je�8Z�K���ADlڨ/CE6�N�X-M�l����f�#7���]0������#��y��o(���\��j��}�|4�g���x/�+��m`�`ŊR���B���63G�'���!�*7p?��Ye+~?�xh��Y�_�-+�m��l��,K�hÿ���y�t�	o��(8��>�p4L\����0W���@��-�T�7���  Bw��lzϦ.��*�E�=��)a#X��:@/����ImTS��ܬۃB1�Z��9%�|�d��5�Ft��A�����P��H�����v�����}0�����q	MPi-�s/�\��'� �)f���ӓl�$-��p"��v��d�)���taK�'�>�o�7�CK�Ē�޶ -ռ�C�l�qK���isFbYY�I���jǕ!X��'�k�$�$��s���h$&��d|��l-��C
�����i����u7
���}�a&��*U�����J!�`���2�s��I�1���l>��������ۅ{QQ�%lmܮ����5���:s����aVkiH=">���LK,;���P��s�!��ߜ�X�57�[9��S��-�S��e޷s�=��6�{|�R���L�3ë72W������V���b&��X��@�O��F+�2�l���{,��� �b_b ��{�/�W��V����.ssM�Thf�Z�~��j�~	\	��?m" ��\�E$�ѕ�_��Ġ����O+�@��DI5�}�h�ƛ�@7P=L
�7�LF���K.z5��Y[a0_h��� D���PX+�(���0�f3��T��U��@2A�k<��xJWeR\t��ƚ���V ���KǷp j��yN&��,ny��dRc(|� ��w���l)�h��b趗?h����r8�(5$�	�/��`N�
�����A���P���a�Ԓ(a1�ڋYG��FZ-��Y�i�G������ �qO=�0.�QE�ZE���uER:���4o��%���j�۠�V�P=��7����i����:ũ�dJ|
�d�"V`G�nt{j��b(R��hdn�H*��R<w|�b0�}�z����q���i��^>����%/d`�p��ٗ�0��E�
e	:|�	�t<�":��LXlxV64EB    fa00    2ac0N����[k��!�H^ ��U�R��=k�
�X@c��v��~x*�B��-�V%
m�0d�Kj����qNr�&و܅�˼I2̣�7lę��R�c�c�ZF�"@����<��*��]����#=��4zXۆ��a�}�am\	��Gu���q�&)������v�Xm���������E�f\ye�K���P�/��wTb�C���Y�'0x���/����+�=��[�L��b� 	����3��@��.����a�c�o"0�rG���5�ˍ��V�;����b"p܊k �T�sZ�ZGˮ�b�N���]�t�
�,�}>�$gr�\���K?��g�e��
	[;u�Ik�L1"������z4P��b��w �٣(Ӈ��IU����d.�ԙ}��Oѷ��C�>,B>-�NX�v�b���)�~n�޾/�k;����(�X�7yG��Zq��JՂU �{O�
� !V��7��^���E3�N2�h�FA�|T�b��2�u/@e�(�-��&z�m��8l�7|����r�+�����7�5vmo�������2{�'ޤ��h3��kZ2��g�	�?'Lb�3�$gĽaA�h]SG�"�~�Y��T8��/������ Zq�_�\מ��T-R[΄0�q�;���>�T�&��i���@B�sY��G��Sh͖�XPNR��l�+z%#ݱ�_đ�s�����)�.;[>�h�CO�C�A���%/��f�
 hw(���nm���X:�5��i���f��� }t-�S����2���=�D���F��aR�����:�p����D��j�xRQ�9E��jZmZ�ݚS �����hc�� ���ZT��9{�#_�x�����o��+�/';`��+^ސ�/㜪z;�r�l�t��{��y1R	e	�a�I�\- n���b�;<���?!|�j�VȆZ��3��ќ7��S	VR����I�JT�_�5T\=R/�2d�����%���)�0c�٫����ԙ�3�2�b����תm�C%{m��
��-bV�!8sR�Je�+��օX����4�࡫�k��J����=W�A5Q�c��B����1��A����y�#:�Kx�ޡ��K������2���FbH$��X<�� ��B�U��[�^7N_�s�z���2����oD���q��(ڊ�4lX�	.p<�8��b��x�Vx׎V�4{�K[�ڊ��~���i7��LzK�e�1�_���<ov�ym6�bA����,T���+�b��Y c ��T�?��
�<�XO�w!�bN���}�;�z/ݘlT�vh�M(�|A䦟�ն=#[r��p@�J�HN^�� ����T���
�@����q�F\���4��t�q��uX-�.���Å55�,uW�ӹ�ĝi`,��	V�����������[��AĜ`C?"a-}5���N�4���)�����Z�TS��.K�x0-��.:�x:ז�7ҽ3��L�y����� ��7T&���PjK>Z���捐����P�����oIu��&>8	���C)?�� <m�z��V}e*M��H�ֿD�(T��ӗ��l�tS�'E�Ǹ{y��5�_|B�o��s������~��e�Y��8즢�v��W������C���Q���`�yS\� �;�T��h��=Ri_W�Rd
�BR��*�_ǮN��EX�A�y�嗊�D�����쫜�A��P"ӻ�,G����	^��'�'�ֳ�HB�c���'��£�?LXf��q�|��C"/D�l�hO���=����������t)���v'Q(�:�h�%B�ܜ�5"��n��f�F�:H(Y(d�,�� -�5A����""�#�Ogv�����=_4�2�R���aoò�n�
�Y:��Lpuxo��.88��I�����
ת.v�?,���W�Hd2.���:��J ���Ŕʃ�!h�`�[b�?�b!3�n�
a+��FB��N��[��ס�: Í��A�&4��s�H����k��\���!w,�IX���]L��'#�;��� =<0~��[b��4�Q�/M��ApE�v�P�K�����������F�28�˫|��{)�1gD��6���Y��)����l�5��~�U��Qy��8���FF����na��� ��|�r�rD��>����p���I��xw��	c����\q����89��:�fM�g�Bz�q����b�H����F=�	�&��ybkP��9�C��{@�
�g}����S�R�6=]��6T$k٩��qq���������G�#g$Gt����O����Y:$J��`k�L�M)(� �V�į#U,\<4j��b�M�b�[;u���J^���߲�����^V�����JLeE^,�Z?:�)�搟]������=~<��!ET�z[�?oM��ln����X���w0v���S�#"�������On#t
�8���L�*�K-,�|�v=�$,���[�ψ�t?��%���Wx������2���o�-��A��*+S,u�v�75�Uw����T����Iq^�W
�a�r{����Mм-�	M��C�H!��Y�赌!�h�tH�E�[��u�E.�`{���B:�T��%���#�:�[̣���ݵ�gǌ���6i�+���:uG:�[���%I�ϡ�{g��ħ+����"R�Y�|�sz�b:��V���8�X�=S���-44+�}�PQK��a�X+=I���by��z\�2���2h�7+��֌��.�d�_��*�M^�o�N��%���9� ��l�Ź�g�M.������R�쁦񙂣Y��Kl8B@Xr�W�:�~�y:��0��]�Ւm1V������,���[��==��e�s�ZEު&���mw?{ᨛ�Q�����W��f����b�v_�cf�=�O&��֒1��Y�?r����9*�۱X���^��)����
���1֦���8��Cq�T���WE����\�p��5�#ɡ��b��b���e%�C�+���@�;�mW!�ATB<�L���S_ӽ����J�!`{�a��5���Sn��|	l��I.�k,�W�8}o#p�-��a�U�&a%��Ƅ/�E�(��/m��k'��9�4��gX���F][����z��r��g��A-9d�-�r&:����,�@���������S��ݑvH�GX!��1�!&����iᨅ��K�>	ƍj�-�-$��j;�	�p�+�g+���x�����_1���CGL�G�1�A�V� �y0Y2����p�ٝ�f4:��;y�����NӤ�0O����n��|����������v]�N	)qh/�XyOBjwGL�B����Ŝ���}<.��90�[L��$�(�J��j������^����!M�\&�RZ9Wp��_���QU�n�h�������v�����0)C׫�r����a����x��]�xw�:�^�rtajޙ�>�g��;�E�g-kkK-j��G�FV�O�j���࠻6X����4DQH�Ëo�c:fW{��Gf� IkG��d�i�g0n|��j_7��@�C�8���:=�������1b�z�	>J�>��ɏ�D�Z%ʎŎ���0W<�Ѕ)nB�j7{����I�h�	uGjNSv�:�F�^�RR�zu�oKS��.'��mx�]E����N�Na�Fг�T#�_X���3j�/-��M_e ?Q�j�e�T���*<�q\��S�U'S����:|��ZM�aZ�9��2춁zG@<h���K���q9pH��� ����dӃ�;ۮ('��Gw��G�t�䦗 �iGZV����U����Ր��-��TR������Y�h� ��"�є�+�P�abw���o���=Ɔ�mn�����p�JB��z��ir1�S��8�w����X$�y]���	Pn�i�y�����^^�`U�=?���X��Y<����ހ��%,�1'�&�����/��t��hɣc�%p
�rЭ[ o�Y�Iq�q,!�FR؛�Y|��UCø�:WRⲨ&3ayS�:SƢh�`|��w�T��:�TDc#�9B�6���' ��h���K�&(
�#�Y)[f�g�2��{w��|��ጌ�ξ[I2�!�>Qs�a�K�d������&�8gWKC�]4}f��IƉR��B��!�7f�ҸJ�{Ш�ݯ!��)�@�Y�H�p!���g��s��hH��d�H=�����D0n�!���u�����Њ�/���㒂�h�I���hgЏ��%{g�u_q�R���a�п��>>��Ge�M�|�Wf���A�L�)G�S��z�m�Y�r� �v������X�_V����Kƕ���q 7�d�ή��d^�zg���\G]�qC��+�h/��'(QdF�#��:�W��B~dfv�cz&<�<�w⛀X�Q�ޓ���]�bUs�V�#vI՛y62fp�>�|��eӎ�X��X�����^Zw��9�#�Eܛ�b)��[]��vķ�CBm���1��qX��j(^�9!x(<��
	ƨq�`,�[���5�������]`�/�"��ۓ큝r�|R5+�|Ki��nf����3�ԓ�.J�%^7�PzMxC���5j����ń[���<sG����Yk����N��:��g�mʴBD��v�fE��ɸ�e})�� �h*�q�Pq@:{��K<�����
�b͗W��ki��rؤ���X��=f�-�w..��E5�g�a�:CrѾ}�m��H��ڧ��f��o����מ�a ]�p��:iA���x�$|�9�2�u�8�E)��lL���⌙P<a���R�:�P(s"8�6��d,�~0?򴇗=�kنK�?�[?+� Hu�@��0�ڌf~�|�x��2�I�����A�M6�&�5M~3-$~tx}f-svA^�l'�RԚ��� �������y�x��K�d�oˮ��0,�Ǎ����2�CƓ3t�����V!I��5Xiܧ��SL]��'�Q͕���������-e��~���ߒ�.\���]k�g��l�5ꡧ�gR8+���G��T	ك�4zDK�o�T�:+0d��ܳ~z���y"F��H��#���D�X!�pg��g��[�n�6f����kCڿ�=n֒!�4-q�N�"0�8ǚ�&��B�����F�W�� �<~ޟd�mjo
0��xg��k�c��	��$�0��# J�E��i� �k�0GZ��S�"�����x�ˠ����B'�z((�_̓�������>���J��
w��w�ߑŞD�z|Q�3
_<�p��{��\ ��c��b�lK#�)av{���1������C��'p�������s�~Q�R◔m� ��0j��wך����2��5�EK�ȏ%ø�J	{hk�4��]E{UC)�w�n�Ɓ :����!�%�%:W䍵�=���K���X�/t�9����T��G��(j�kyv/�:�a��NN���SFˀ�{�iu���|�kH&
-�%���z�
q\���v���Z4�ݙ�xu���s��ZF�}�4�yOO����?vK��?G*�ֶx��� �>�����b�>o뗒-P���^�0�x�6�[/gS�g�
躛���}_�o��
�[?J�N��&��`=��>�o|-����.��v)[J��	����'S��*P��=A5���~j�N�\/Ls�FI/9���̅��{[{����I)B�%*�ۮӔ(�B�F<����H��PoXy�Ċ�(1������jӬ�CQ�vj�����5%r��L$p��[LRS�4����g�ضTm��Wܿb���a� a���MќP�v�F ioA ��8��݊�}�r�����*d�L�g��ؔ��P~m����ēI �t�����(H���L9c�*����=d��e�Yb��`�c]�L���q�H�E��0�ՒF�������4���#h�d8�.�Pi��,����*�G�L]�Կi=]] jh.\�����2�S����+�,8�r|��b���&)��+�7I{�5P�d}��.e��R�#$�	�a��g���^4�C�|I`'0<^>Bas~X}:�T@-��>�������%&&�l���C���AK�稥����r��UPv��Ұ�[�E[e�{B/n�ͮa1�N���R����� @��yq
(���Lgx���T�嵂�cNb����&?ˋ�*nE8��[(�zz�Bj��v�� *n��c����T�ɿj1�7���lqlĚ�R��Ԅt�mn�}�xx�����EH߲ԹCN;���ڀ	.�e�fu'���b�ὺ��J� ����tr��U�b�(W�.w�d	\�:��v��0���SP*�����W�ر��<��\�'0g#,5���G�����4(�DG�OP}M�i����.
�8	����V���ʧ�Ҟ����	�	���!D�{:�%�qpx ��4`$-.�Жgs�7b��Ƕg�e��V+��Bs���s��OT�sfu��7n�H�}�1A�w�㛭���lG�iP�z�eb"N>�.ʑ��}z7�͸��vg������� �y�#޽�peʘl�H@"��@�^	,Iv�� k����IF�y���e\b̸�����Y
�qh��cx��9V���&���x3�2��8
�.��WU�ܦ�v=�w}���|\d,���|W�B���m�@|V)���B���:ɘ��K),��f��+"M�2D`�ޅ�@�#(�jq,��W����9W:s0m����G$�t�3$�A.rS�~^L��gK5���$��$Eu���&oמ�/\���b���a�z�A����v2k5��@z���z�O̖�.v6��^Z��2J�8������Aψ�'A�D�B�G�V*4�UO���z�z�qC�e�h�{Q�d�O���o���7~z�P��A�u�f�`�K�@����M@����d�V�U2���|�	T�����,��� �s�i@7�d0�f����R�3�5F�h�A��-T��P�d4�1�X��H<`�E�(H�&�O����lKۺѫ<�r�l�v���y����n ��&F������9"L�{3#T�u�V	r<���Rz�,5��Ck�2�]�њ�uryw�<����q@��d�K:��S�Ey,Ң�:�ڠ��^k�G��,���[h|>F�B����8������ť���V"}�\��tU�4�.��{��TN�]��W�A�xhT<ԕUq�Ͻ7(�2#��?�>�G���&6r���K�ca���G�����M}f�_���)���� ��|�Z���6�2������V��rĲC��?�oj�5<n*cSU`whI�@ �.�����b��7�%��H��S
��=�"6U�v5߃,�.N`N�9.�\p�����w�F�X���s
�S-�T��(����`�Z���Z9�?/R�pb��8�,�Z��p�����C�C��%I�DU�K�B9��F�K�cc^�ղfÈe�`�x��������;���*�=u]&���U{�܁F�L�Ri���P��x w�y�?��b�Y�"Sن���pj��05	�,��*��W�0�<��O�ܡ���	�[�/a1`A�^�`���K����6\]�}O�"96��a>��*��S5�~�\��`�;�q>2����S~�	�p#�����8E�ީ��et�2��k���p$O� ��,�u�9���rX@�mwE0̲-&���\��x&Oļ�B?�vp�s�����iB�k��5�=%؉z�B� �@��Nl�=��� ��
�XpN�����tߠ>9$,�N��#+a��f���}�5�<h*C�5`Z��`\������B#�;;<8�>��"��������鷣�.��6�y��]+���*��9�߯�*J�����Ow��������.}A��}b�P���!��N�KH_�7�9�=�Z��EWC�W��N<� ᒈL��.�ꏔ�~n���b��7Wm��	s=�Ҵ����.ˋ
2�#���qC���cLd��5���3;�݅>��b�sٗ�vp1�8�����(��������Yp�l�JAgdKX��KR���{�qQ3�#����t\-@�L�Jc�T�ﵰ�(f`S1��(�v���A����QQ1��]r7���r�K �������"%�+K2���?f4)0��6H´�W�|G�9m��g�I Ȏ��E�|��Vdf���pU��Y�Y������d%��!އ'� ֈ)GAuKəF)�|�44���JK�%��:
m1�˜������2�Jb��u/�)5Xߝ8��cIjUz30�E�,6�y=*���iNSG���B�x�����T�Ǵ����6/wc�r�ף�
IL�����Y8#��������_��K>jTs�%�S �B"H#	�I�mЈ��n�N㞨��R�+$��X���?�=�誜�ƣ0�x~��R�"�oNVC��&��?�;50��â!ݿ�>�mԇ���<Ѵ��.{#����W��=��)틯��-S3�=���)2E�Go�p!�-`o�*f�9\��S68�U��Y�LV��F)=`\��՝��|��R�������-���V��X�p�#[n|�dn��$�D������2|�Oe��0�@<d�UBƞ2�e	�̇��lڡe���{p�x|n'���2� j U�fĸ��8�G�v��,����r�Ro��K�<[����Z�`I�<�d�3�kP�˄7^Ҿ���n�:.P������R����А.<ʂ^<�6�� �HW��$~:��c.]˕\�|���-c��E��44��0)��	�ո�2�	@Z��Ɩ砾�A	�~k-w{6
��csxNV^�nA����Ƥۗ@�9���@��b�?a�ĢxS;��+C��9��tW|���7�����a��ǤHy�>~SY!�2��1X�����A�o��#�2��a��v^�<"�3ӈ�?���{N�Z������u����h����gNk�c�Ŷ��8W�j��EiY���F��H��ְ  �߬\wz����Έ_=�	���������>�������:�&�3e��xل*����\6W���	n?A�U��ۑzc��
DB �`2�j��	���E��;ـ&�"��`�_<v~���D��<	�wE%�u�>.ť��)��3a����Ze�O<���@|}��p=�5����`�xSg�Q7�Y��4+>�u�^�<��6P�y}��#�!����5fU��sJ�ߕ���5�f�ہz���p.@�d��/��� !o1��d%�C�zT��K�*j|��,ĭ,�/D���.�L�pe�N�*r3 ;�J��um��dL�����M/�U:J�\�I�+��ݫ�R�yr���ҹ��|��w9{R�?��F�?s����=��ϕ���$��B�&�(�ba��>  �Ұ$�s|8��aC᮰w���;�7��r&�:,�f� �h�����Y &�B��@hO}ox1`)���`�+-r�Xy�6%k���]������<�{;M���7� �Et���z H�n0�����]]�=/i�~�0\:B��b���E�q�(FWޘҙ]���kߘ��ȪY4kÂ1;��m]����}V�"5��������O�
(.2��C��>c3WJ�Y0ޞ�rф�Y�PZF�����X�S��e� g�VڻA��V���\h�ˣa�_a ���&E��@?��D��bX��v]��4����͂�����\��+�V���_��,nvE�����0!��o�Y���D��ak�>�Fkx�+m]@��T�:v�yG�2�nz�lr�	����#���H��%k�*�.u��F6��fF,��3�Q�SU��ڛ �M��}y�ۚ�� ��#��d& �������	�]������J��^8㇢F�f+1�&��T?�lcbi"NjH2`(Fx,�<�v3nv.���"y�|SF�5W}�GV��d*���;��v��� �?Wi+�99e.��S����tv|n�y>m��*�ߘ�Y`}�h��BJ�?w��g� :����\'��I:y��Ĥ�sk�o���`��}�Ė�=��HGy����A��g���эBd�?�j/yT���'\�1�rkaқ��t@u�O����{����-/]<��3���-m�ǀ"2E���jF��#��.�>��z���-�&���#���"r������pk���3�.@2�[q1S�~=�-��1�����Y���N?��kS�s���ڌ��%ˎ҈�+n�i.5ޚ�e�7�Ԙ�դܪ0c��Z�;8�tn�P� ?�w�4�*����% 9�R��>7 �����V�Ґ���ڸ���n�k��^��
����%�R�4�yPZ�����g��u3�-�'���-����^qo�?+�U�K����a�CP\C�U��I&t&ϴ%�O`�C��QN.�234S���Q�FZ���S��bC�o0��Hn��pga�cY���O ��	h����,?�8��h�z�=���f��)N�f�g��=�ſl?J��pd�12����i|��5-�K	a^h*,G�tjsJ�f=��Q��6.��B�E�?��3k��S��ndc��7�)��=�'S�����Lf��Q0��Wb� ���n @�KI�e�8�G/�3��F�2t�,�0P;o($������w���������Ӟ����X_�� ��m�uN=+H���
���@Q���v�B-�����XlxV64EB    fa00    2740��5K�r:p�J�:�0�0�-	vFʑ�
��l�HD�x�g�l�_p�u�>.�����sh�~"Jz��u�}���h�j�3������Pz�R^*�?Vv�!nR���������,��ۺ6Sӱ����x!�,�h��>S�z	i�4�ٵ��zk�����vħ���g��`<7����xͲ��%���Cߠ��B�m�{�����t�SCc6�8Q��$�#��j�R"ӻ��F���x)��Se9a�*�K�,
��������3lp�,����+͏�"`�����S��{w3����y���
>��y�|&�j&O����B�I�f�P$��f7T��	RM��2yW������!�Ug�z3�ZO����-l����j�^u	�MN����oz���ec������xL�``�7fi�)��s�?o-0p��?o1h�*���Fd�:H�9�d�c�"T��u6�	R�.2�gX1I&xH
_�a�ȩ3b�L���0�����1�s>|�ҟ���'�[�e}����>Y�T�<�,�X���_���F,J���Wu�%�^��G/��$�E���=a��� �WJ"UP��5�^���ר,��W�Ӯ�s��"(ꃘ n� 3*�[�TG)��Fo��>�L���u��>�@[�r�32�ѣ�/O_��u|��5;����5���bÌ*�&���a�����[B|�>��^M�Kp{�<%`��Nq[\U\ #FZ6ir;>]�[���D��}�D��hч�O�'����egY4�)�d���8ϵ��;	�*?4?.T"H34�I:LL&�z/g��2�8!�h�:�!�;��x8��0N�gwp�*���]nl"
�.�Lo+�p�W1�xR}IC��9p �b�Ö�}��J�*���Ǉ��������\�����&O	��W�gZhQ�j�� y�)�4YG���;[l��L��vdu��v�/��z$�h���C�|�2��:��L�P�[�}A*���v��-8�ϒ)A؛�`!ZJF"8j�t�6/C�rp'�&^�$p�[�Đ�_\�!�X��:�� E�
��Y���ё�ßßLa.T}�v��Mu��R�R9�p����Ե��a���Qy�&��@�q�ew;d��	�S%/pg�3:��HT`�f�����:��Uf���6��[b�ܥ�tvYL2�ks��Ȓe�)��hXb�\,���H�Ǯ3�-q͆6��?á�s���;��i�E�I>+v�ic��d��LĨu�Yjw�!(Z%ȸF)Qs�󂄻���1y���H�� '��,�(�����H|���	�A�Д��L�Ƙ�FXM*fjjf����Do3�E$����4�sS�qg�Q$Rk��|�3������M�}=�]u��s�I�&�bb���m���I2�q1�(�t�1�)o�<&g���O�h����*��p���2���7ŷ�k-*5���+���Ydhq˰Ox�w��4�#r�%0>b���sE�S�}���2�Ԓ�R�@��}��!XQ*�l�Q?ߑh��#J`'d�(m�Z(�"�	Ol���Z��B�c����K%|���'\��pZ2 ��Վ�R����RfwN`�>k����CQ��.r��}��z�͒<��%-�A [|+vC��yQ��)1r6Nn��E��?>@Yd�|.d��ߵY���[�F�Z��w�LXMc�\���3�^���x���8f.(/OB��+�2�Ӱ<�<sQ�yX�#�BoY	Ғ����Rw���5�p�2��b5ȷ>��Ь�Y���^�ѱ�1e^d\���_��U�}d��T���3�������_�w���͞)G��-�d�����6v��mX� ��`�y{�>zS�;�����z�V�5�iwY��� �x�ʮ�w�ޯ��o^!�A�K�/�ד8�뺩�z���Br�[��V'{���&OT�-�j
���	�'������a ���Oɴ�W̄��%t'�|�	���d���h�e|0|���������n������{����?_�Ҡ�K���"�g ,��!��ω��l�3Ӻ�Z���?1���Ç�ɟ�Q/�1J �	7�?bn�o�i�W� �#E�������j�(�]Bj�����,n�y�1&uh�Ac��� ��#^~;�ъ����ju��M(v���mQ���J��@y��$��!|����`�'m����:\���_��k)CF;��M��Ey������,��PQشm"��� p���J%�����)� �M�G����>ܤk�M��H��V�q�QAbJ,O!F
�W�b{�bDe�P�	�c��)a6�Yk$�dɣI�x>Xy�I[ܽ"X�P����'�5W���w�Y�J�j�>ײH/�
a��`kıS�F��������!��遫��.y�ը��5� �������=u�@'��_�!��F�g�du�n���ق_~9�a�v2�@e�xa}9C�U�<�/� �O}d�c)v��b��*g�&7.N�q��t��LR@X���74)��y�JLG��p��u�?0;cS��r��ً$cy��`�?��Wz���=z�HCb��,��j�c��1:���
���7��~��p����{8\�cI���k�۬� �N%�ZH�[��|��I-O��Ze�T��G���� \>	4MԆ6nav��,?�9�|@�0�Ss�Jly�`�O�d �m�	�(Kw��o�S�n�];��=C0Y��t_�	g\f�a�"��Dr$~�٨�2[^���Ec�Vh�xzk�?W7�<H��wgW����g��h��WO�C�ψ�`f���ѵf �׳�'�������N��UR/:��F���\�N�M�&T.&5��W����^`Y��7N�yۥ�nq��b�����d��\���/1����W=	�k�/�����bFx����g�m�k3�������mkszkzՕ������`��]��%OG�\��5�y��/�*�Hf�0u.w��k��<K�̴���q0�V֧�w��g�9�Ǚ�����@�|̷U �;�Vk�/"�{{��	.ueD���k0���T��	@zT�?�6���I>G-2d&@j* �o��F�G@�'�D��V$�ZC��|t*l�9/e�|��^96��Z�In�έ����kB���}Rc��L%iT��=>���By)�Ս/E4��C�������I��vF�`Tb�&�R�n��x2�NC��JT��V����T����
Q�CN��8Hh��̀���W�L ��B���_�(�
�A��Y�T�Q,��/Y���9�	�5gEr%n�cy�IS��x�B@qs����{УΥ$e��4�a��%o+�t�1�'y�E�OCi{U�0GT��`8���Bsp� ���C���>�:A�>����2(7���LC+ByFs��-.�D�ߓ�c�Ƙd!�T����2Z���)J�'��Et��i�s�7z��^EbKA�L� �B@KWqx�h��4!)R�D�/fR��Rr�~�����dC$��Z��}���c䁋�"�����C����l�K3�ɟ]�rY��Žn�):gT���r6��ƒ�.䤉�$�Uŋ�Z���������Q<� �U}��KsW逋��Va�i�l�g��f�2���/����ʀ�e�紉�	���`6!g����`O���ΰ��.��C"D�䕻�뻿�'J�a%��&3�����I�������a*�r�\�8�(a�迧n	w��-��[/��M���Kw%�I\zq��7�2�=A��D����Pc���s��P��-�4�dX�3�n��2�w�j	Ly���eE�/�|	�-8i��Ka9����Aǜ�wuJ�
���|���KVjf���`2�d�cm�":���@��?�b'=��sQoV�Gg����jDK:��{�+�|RQ����,k���D��,��8�]�R�H3L�CK"�3��&)��|� �����~��#����Gz�V�J�z���ȔnNGJe���W�X�I�Y��	E|+x͗!e�
iS�H�~�T�W���r��`Om��b����-�
�N�|���V���5��ᜅ�P37W&�#���Az�M��:|�4f�jj@�M��̹=�T���H`��E�����*<�l[^��z(X��f�퇴X�����4��Qi!jqu�����1�$��t���!dqj�u�X�k�ݹ��1j����t@��nH����y������؃g�X��AE7�X~|�A�KSXhb��yu�c˨���=^H���YqqJ?{[R���Xwk*V��Z���I�TmiWn2r�{*�N#��T��G�+� ``���fL_v�·d��Cȭ{z���r�2���ẁ�E���h
�^�N?����j�3:�1���x[�{�:<�yϤ�X������2�]�����!�6�V��R6!�ǲmQf]:'l� �]�Fp�,E)��
N���;�>G�J���cgk��	g���U$�R�+/B=T�(S�^IbUv0����B.wVĥ��ե45��-2*�H�x&����N��<��l�DgW|[�͋מz��B����UP5nyA3z����S����+*:H?=#���e䞳�Y��
����07a�k�,jS�����}�v�o4)h�����U)C1�yh�����%��j@V���(8�9��A��	�������3�Sy[���yb.?��Yc|�D��[U�t��N\�8	UW=�1ԞZT��z�1d��v��P��и�� ^���&r�>W�� ���-���D�5��P5@���7ݧ#��ƥ���LZ��:���-;_�Hfi��8yh0��&H��'�d4zA;�-d�SK��~�dw���Yaє0�0ԩ�|����z��wܚܲ�+Q�p�^΋�v��$�f���,�������G�mD�ڟ�s�Z#�J)`��)?B����(��;��N�����ވ��c4e?�����Y
R�4^�L/�R=}"Ra���'�}�m�_�qtF_�?��Zѵ�.�V3�y�[�3���^��<�0"6�g"id�j�[n�l�$'�g{/
�؟%,�J�q���p�7}��I��[��b���n ��B��Ar��XF��'��V�a�H�G�����[�ֆ�t~���S�U��%B!6��Q�Zm-�5��lRA��� ���
��Eg�F�H$��!���t��S$t�]�2����c^c\��$5E��^��l�\3FaT��i��:&a��I�l���ڂZ����bS�s��y�~A#-�l	��q"��R#D����ޱ����4�ϛ}{�ПIƮbC+*3`������H|��+Ǉ�'�onŲ0����	���O�޹��H��=�(�Ke��#Ԣ!Ī�=�6k8����Ҳ�?7A�=o��00�U�q�U`D;��F��}��M�YE��`���Y�g���[�������6�VV��ȋ��*�UHT��I�7�ԝW����6r��<��a���:��h��Ɣ:�F�sd�"�fi&Ԙ��C��J���73�<�X+�-gkzb?7��,�q���{"����&����p����u�E�?�@��S�ު8a\VbV��1����E�X2�ᰜ�(T�o/K<�ˇޞ�4�pO���9:e��ku�4��	ᓜi��y�^�8���+X��D��@���L�+w��q�J��r�G��1a�!���T��T�ۮ�`���pc՛o5�Jӭ%�N��,��A�s��ľ����o&$�역g�HX��/��!�0i_��_R�KI��ƬR�b��}�4����?[��輟�".�����-���qpq"�sW%�7��5D�VA��ߑ�
�8�s5=]�j߿�s��4�ҫ�:��8k����@��~޸1�x��&	a��Z�$����k2=k�jM��]D'+��`�~��I�=N���l�O"� �nT�)6M��K�D�#L�;�D��z���ݶ�I�Q]�k7����3��Õ����̣�Pm�[=g��CzP����	+$(hF`FϚ!Q�ͫ�@�զt�̠>�p�h�i�T?�DW�D��� �N��\��=�&�Qi'�%��	�F��*a|���bJ�	�����,���2�[�0)}���)4�ti�4R#�k�rfQ�muN��o4SE,�6�;��,�X.y����fc��D���f�+'�i��7�+�f��w�g[_��'��iΣ���Q+ڌ�xbPdD��dE�,w��t{�s'�Y�1�̸����戀Ly�m�'*=b'm��\oT��u���ڠ���U�>�1�`Q�!��݀o?�.*�P^���s���-vN�C>�[�c�A�iE;G��b$RX*FѲ5�����pC���^�]2X (�^kl|^pП@�}i������%��ڋ��d濃p��.�`S!��\Y��0o�6ѻ@GT[��ђ�t��K���u�
��A���5	z�b`��m�<��V��U"����32EJ@'(�vV�5�/l֘HIY��^������׳5TZ[e��zf%4x�G~�v�����h�"^)D��n��wtV{rY�t1����~�hoٷr��՗UGumȍ�R�YCC�Y	�7)����@7}{2��`�+��W�3��m�W���1�bߊ[��;�2�c=X���׿S9��#&��F>P�:!�`E�PS�Z���Mq����nkiz,��dphY|�##T�����ڶ�Şv��,=��� �bU�fl"�4]+���[�#��#;��^�g50�)�OM�*��:�3��zW�Q���%��L���iuB8�"��~�<%*����:U�<dFS�n�*C�$�:^-��)m��f/�{'o�=�F�sH��/_��Sٶ�'bj���or�k(��ҧZ���e��Y�=�m�G&	v-K�Q�ዬ��5��B��+?/<Z�!v��t sq���<���E<M�!�nhou���Vl��Z�BJi���#���C��
'_`_b^���D_]R��@�wͦ�����R7+=�k<O8��i?!n��V��]P뢼��Y'.�ߴ�j���L��#k��B��0�}k��=iF�e�銣�9�<]D� �����u���hz%Z鳨������ckO�:_�r���/1c��P>��'�(үZ�t�r�lA��j^������Y���H������]M�H|��j�9_����a{"�i����T�>4�ʾ�R�����@(�9��|�PE:��d�D�*�8�[~�6ߧ�"Y��T�b-$�:��k\��~��<yd�ٮl�q)~��Ʋ��13���2�s��]�����G'���a �����cz���
Q�
��4;�id���p�}��A�/��&�oYJ����>��S[��}�ɂ���7UzK��A�.}=htF<�'�u�ܽ֌l$��gJ��t,��!�H٣��8�:Yz^m�|��
A�H�{�6��p�6�/�hm�Q�U�#^�!q������m���8E�5�	��H�y�ˊ����!D.��zą ��NKl(/0Ŗ\�&���q�t%�+�8;�����x2x�� ,6/�����40�,�?����W���tS�"�ڴo�䳠�J����<��
��u����>ͤ�����R�@'tܸCs����js|�� ]]�ѻ{����X]�`щ�����K�I�K�i�<��+�XDi�qpHiK�?�eú!F�Jea|G����hH��Z�GZ?o(ăN�AL�%W1w�܎�}�6�R%(�;eצ?����E��r��\1��<9���b�J+�j���v��|��0_���m�^�u�3D^y�0 �z ڬ�2S�g� �Em�~3pE�KɆ���f� ܩܤ\�v�O�޽;�J��cL�~�ƍ��1�4U�	��H�O��NjY���R±bn�ƻ�]T�F	�=��7Jo�r�Mz��6z�&�~u���D�֊���u���Tu5���DH�b�ȁ�lxhj|o�[<��<K�q���8��d�v#W���z}�����5�In�d@a���[������U�|���g ��"��[t�����u�����E���⢦E ˔�3�})g�w/q�/���ߴ����z`]��൏��1��]��`��2� �.�NW�0]aL�A���L�,4S&,>���^�G��^��-����
��KM:P��	��+L��p~"|��]�3l�%�͙�#�!���*l7�x���"Z��71�h{N�mB1�C��^~�e����qplsVm���ɔ%�ݩN�v5��O�,Ə*���w��
Ce~#6���cc��o����Z/�ϫ70�W5镔ɦ�"��ħo��vh�t�=M~�oZ�uu%��Y{�q�����'�?����6�t���ïny%��E�:?nou�C�ne����v���ԅ2�1�Ns�+�n�~��hj�`�c�	�*V��(>���L�Z R~k��<����P�6/c�7R�'7>���NTѿ������n�s2>���e��C�;8ά�a�ƾwM};����wG���Nq�7v#�q멑�ݤ�P	�5	#9�S���f�M*����x��'I�1���m�J���K*�����U�,�:mŸB������r3x��1�hS8�����(�u����"��LV���o?K �)�Ȓ��K��c�S2 a���x�栉¿{+/E�8ˉ� kG�oA���3�J�}Y�c�e���t�a��++��:���2A���pv���_ax�_~�9�C4Ƭ�#�>�ȥ��nV�V>���Q�+z�����:QF�[�����= qf!n'VNG�����"w
��k���>�Q	N��������u�YX�Z����J� Ң�4���z��A̪������G�L�w�w�׏�=��a���;��^A	f.)�=�tL��uʗyma?�?��A�MDC��M%l�V���m/�����V�^������,���҆������)�q��ݛ7�s0@�,Q�?S�����v���P�_e�j�}n����_����G}؉*��	D�nri����Qt��Cʭ��l#�g'A%�Ւ-�W|�e�������d�7�$����cl�H�6�OU��*M�~�$�����l?]WMB���� !Zā�E�i��U��/�Z醾������vU�DY.wO�?AaT�C5�������;���B�	�aB@�EE����qg�>ΖW��4�mU���J�� %ǔ��W��:��j�H�C�<f���x5���o1~&O'e�����9Wj��-���I@ŪX
��s������v��^�(V�χ$9x�$��lPR?��FweN�#�J�s�J����場%�O핶��+�Վ�2����DbEzJw�ݬ���'�8e�3|X������A8�*����G>���t8�X��Q?	�i)��=��3�0h0�� Ą!��\�~���Q뺤�7q��r�	��� �I}�8�zK	YFnۭ��zETq�y�L2���0����/1�$w�`暝��)ߙzZ�"/T� �y�����:I�Lq�H�k��U�F��K�sη���wKޮ�p]LS_��.�F�I����
���4�g@E1u�w��C48��5Q�d��+�mL�ra���~����w��h&U�R���ڬ������I�����O5R�*/��S���rxU�.4��6a������f����K���Z�'.DrQ�~pZ�W�LA��I�����a��O!�����Y~����t��?�k<�k� �����&E�7�3�>-m��ZM��`��L﷼�)7XlxV64EB    fa00    23c0Q����'vMb��E�Ǩy���c�,�alg����W�Ÿ�J\2ڿ!�+��4��Gz�AGK� ��r��\A���|�F!��	��#X��*�o���)�߅�Qj-�E1�)G��1�O���dȼJ.q�:(3!R��[�=}�6�Чܘ��V��F�X��pr�i�ƽ��%��e��*���	�2� Q[
7���B�,���Q���96HI�-Wh�3L�����Mz@�xP4��`Ӫr\bU�=� �)��۩Q�*�f�-<ܺ����h�_��?����Oe0�E�G���^���q�:�{[�۽��2����� �?_�T@ͤ�1�qͭ��&w$��	�O`!i�;���\��lf���R��Q���fa�0�/�h�i<4�.UoXP������;$D��_� Y?���8��\�+wq&�q���~j�+ĄG���ѣ�2,��]n��P Qn�a8�Hi�&��AJ8B9O�"_/�7�F�WRudGܻ�9�]g�*٪�|��������q�����to�([~��D�%IL	���;�E\��	NBv��w�o��N�ʑ8�eI�w�?b�E����z��Ry��|�'������)��"F�0~*���r�y��yũ��C��3�����lVC�U7p�i99���݆ts���J��Bg�J���bQ���6Ф��hN�S�C��M��	��ëMg �V�Y/r����Am�>T2-<!�(�1ёK�dtO�>zq?z��U���7R2�kiۖ�:��a���Q����2;y"��1�F�Fg=��'bp�{���i�g�,!W��L΢�P���Wڃ��Q�B}�{���U�%��>ʎ��+Z,��T�(U��Zù��yEa۠��]�s��
 ��#�Q�
8ۡTi�p�d�������^�)9�HH՗��PRB������5�����k�^��*�
v�'��;��j�Ya����鸮��zm����-����L��r�3&|��b|㞍�H�����֛�b3~;�/ӛ4��;��:��\��"�b�Baڭ��n��dL��}�".����c3�*}e����w�p��Q9-ӡ�����0<��������/j^�l�&ָ)��o^�`"���~�;9d�w�����f��R4�B�|��2��%�yU� �%l�v���؟�M{3����	���Hd�׋}��.�]��>�i[�4��WfL��t�H*|iP �<b�!yU���r�\���Ԋ�n��!�
�m�G��Vr���[e^I4=����5?V��>!9T^IS�F� �E�}j��
�[Gu^g}VO�xp�ؠ�^\D�F��v	�����8����,�6Ga����:t�;�G�SS��ڗ��H9!����
N�?��;�`��
���[釗��QqLPm�5I�Y�;�pƋ�-7	�v#��TYb�%%�-�ԑ�?Kb�G��kg_�D�;�j����v��\�h�ѫ�q� �/y	 Ǭ!��@�GW	���.�Ւ�h,.m��3����#:���z�P�'�&uܢ��Ks�&���D\�e�Vi�Ɣ�G=�_����>E_�-ᇞ%m
���G���6�� BU��&�9��Qi�?>$�^��o��!�G���6�&��(���Ao�n�ƙlbn�g�_�v��.��&uz8曖� �(;	��S�E�Ɇ����Z��	t~��k��W�|����5�b��uY E��M�мE�v�v��fql
2?�}`�@���$ٍ��_O�si8o�-�R��EA̟Q��$9Tꟑ��ތB��}ؼ�u��=4�U�)g�?�Nt��gJ{�I�����z��ұ����H���l�3E��a�r��l�������Nۢr.��&�4�L�����G
�:)H�ye-�f{q�X�����p&~]�ԚZc<�����m���Td�7�XZ��;y�.�'��t���|�}�2��\�O'`�=�����?��>a��+��oĴ�D�djD}ik돎�U�n���\k�RtU��(�+� :���Ynt��y�fUB�������^	���*D�����s��hz��f.�.�vI��H-*�[uM���R�`E싕b���HJ�W�3�߽f�F��`�S�P�
8����e�B/�H�.Erim~��lY�!�2ǟ�!�R���l	���l��v��&��o��_�g��3�74OcpI��Cd4O�n��E���������Kk�Æ@� i?�(s7[�k�����3�h���������C%��Il|<qC��� "њ�Xr���N^/�I!��e~{�/`�ʆ:z��b8�G���$g�]0�_�m$Ǩ4I-��ft����^p(~���ꦍ��^ �$錋Q�>�m��|>8c�W�y�1=�ַڪ���(f��N��K!N�*�����Bd�>�e��b\r�|��e�.���n����`C���v�]��񞅢~��|���s/��pv��0x�\���C���o�B�圈4!�P�L�TR>��0�܂���y�W�<m�_�U�
�Z�����U����@-�N��h�S����n�\a\	@?��mPQ����{�d��\��#ި�UsT`���&���%{�V�Ԅ>��H3C�W7��]=p+��#6��=�F�$2��S�KR�U�����|���򥣷�^�~�|�u���3�,�IW���ՂH�7va����e.�N~bx�7xW�-e�bH=�����tI��Z�a̧A��pXܷ>}�_��na��r����6c/漟2�����'�P��42fʫH�P_&ڤ1�>A�^�F���@b�PFJ�?f���\��kl����v ������K�mzo�#`�S��q,�$���k��|ǩ]��@6J�xg@%z��]� 1�OÓ�2ԮZ���Ǆ�9�C��-cy��Vn+�ḑ^Z.9�$��m��QK)/�.��{Zh|�Ϙ�,����U�ګ�&�����H@@�j|sH�*x��P�?&D!*�s�{�pct0Z��n�48s����9�J�ꎪ�Yr3�Y���'�l�>���C����Hn������_Zvc,}���D��P YMG:���@���ۯ`Iqf���8y�H�_�0YYk�������f~�,��	��6Yqw�
�s�æ���]�WS�ޫάXr�@�-s��tR����h�\
T3����Ɲ� ��`��U�%��P=jz����2��賶X4
�dw�`�Q6�9I��ɖ�C�M������!��O��pF�'F��f���.����t~��<C��{dt�2��� �D"$�o,�B���@����~;_�>���)�3M�Pۂ�C�.��{��ڨi�X�Q��~�D:~�,zNICݒP�9�Η��W�a+9z̔��5�$Q��J��񤻭��T~rN�B���i�F��	&Gt͵|����i����Gw<�Sj{�-���܀��0��
��1���w��Sk�ޕJ�6}� o��5P���yN�+�q�;�$N]7�������~�RެG+}��t��(mV�[	��"�Lc�^|:�O���#tiT����rp	-���4=]�T�?.�566�J�R�����4&�ٗ�j@β�V7d�@��Wx�3�oJ�[�EiCE����TZ5���&�R�˽6�g>�T^�5��L�FB�HM�w-���e
U��0D��u㾉&!�n5ޘ���7�)w���X�՞�[{z-��>Tp�4��c�e<;�ۆ��
��mLyq��LNB�7�i�������{;��n�fdYv���@��]�nV�q-��eKV��)����3���d��]u�CC1��v�g����0����{�y�o��{E�"�C���X�q>A��Pޙ����W��`�hMdI-���5[]7���\hI�|b�`�.Vd�+S`�̪�F�(�\����E� �ɇ���)Ni�E�J��0q>߄�8�����ɕi�R����&�ҞꄽP�>tٵ�Dd��2Pѫ�ܗ�W�4MwF�K}�i���>HǣL�G"����ܗ/ݞ[����O��&��8���U�^R�3��#B7l����!�}�g�5��c0	�:A��f�s��-��H(�/=��aA�_�Wj�&o�p�ȏ=Q*qb�n��q��[q�����[�7Zb)�sm!�o��D�M�L��"�B�s�� ����sΑ�~�Z��~�h�7z�y��a趩����$2a�u� �Jϒļwa[aT$O}*;���H�vQ[n�}�Mj⫚K7;=U���Hq��B�i��2�t�|�fN�6�C�n�Ds$
�B߿ Z��^ջ�q�2��987�c�z,�/�݆ߚ�N��>�9&���{�de���I5f42���0�\[oQ{۽���@�ā�oV3�kW�5�*8~x���5&�&�5���⦍�t��n6��{�>�xhMDU�y�Z�fa��L�|I�'0�q�4L�@�k��g/*�=Oq[�*G�@����-�����5���R?�J�T��T��aNɭ��ؖf�s$L�BY%����`��Z�`
�ñ���x�)g0&i���Ů��Q�8�]c�]�n7q�a �Цe�k���z�h{ơt�����#P��j�X;|�����,��,ܓ���g�r.푴��,����'Hk�&G.n�uj� o@y򊳣��nGU3\IU��L��-��9ʽ�3����x[B18�I.���<���k�0I�����W�K{+c&���h �"�2G��<6(��E����L����p)_�m"x[���0J�~R��d	Y�������f�A�}J�^9u�(�a�'I�9z^�6���!"n�,U�����Z���j��Ց�M_�k�G�;�筐�9-��qJ{]{;�*���4����LIIL?����E�>0����SGy>�u�в1#��ݨ]�6���l�sm@�>h�*�3Q0IE�u% �ت���
�3���m#�M�&)�־�3F�o;7�A���$ЋH�� !�����݉hFw^ȏ�Z�ܠV�fh6����r	�VA˙VK����օ~@��W5�N�w��Azp�M_�.ݦ�;�~���O��4�
�SWvAF���yt|�b�����^X
,֬���t��8j�5˚���{<��/%�|j�8���,�
�BłA�&�c�{������6�zrsp��!
u�ٺ�5:�0��46����&�CrĈ.wc$���r����e�;��1wi�%'qK%�Gϼ�j��Mo��0n^:�sɐ4�㶺8�옜;6]�P_�^�Ǘ�8���#!�,�I`�)����)��B2�(��X/�X��*��4��L(\�T��Qk�� ���Mb1s�IR���+��/ãT��ФޮD��'��:�.]����d	%��m�?i�2+S�->��rY�Qw�5�ۄ8Ɠ�X��ٮ�����+K�с�O㓰��.��&����mA�I��B�����@)�@�P�Q��TŬ��7yB��a���9�NY-F!E`dْ_U@��l��?X.��b��4S��a��K}�=�"�6�キiZh�_��Toׇ�(�d�9Bگ$����@��N������^����fCn�$�mA������ٽG �@���J7�j<�����S\Z����Ս�LPp;{�X��ّL���@��NTp�x�A�dR$�� ��oMdr���أ&�j�w���~����F���DHʟ���������V�|}2oZm�#4s�I���� B��u;���=��ߙ����ؚS�N X�,�r0��*�23O#x�lH�L�0�1[�
_�/"��^W�R���7L�,<� `������'�<����Op�ʥ�Qe���c`��)��� ��aB#�[	����h�)CH彂��'���6�����n/R��Z0!q���"X��ϩ)���<����I_�(=��i3���e���3g�ɻ��W�C�S�u���Q���wx�8F8eу�i�|8����헓n$�0ٖ�U�eʈ82`��(������ǭ�����p�z�tE��_?�����"�`v$5��C9B���fN��XI^A�	�h�@�v�޳����X���c���mA�����U�8>�I���G���~����"@'c�Ŵ��i򎟚�(ڏ�]&Z�%��]�6X3� �0c��޿ �=�e,T���:�^Q�n�ᑺ[؂�,���Bi�a���MhHԛed��ǥp�,���b�����R�Pu$��� G����ܙF��r,���: �C�̯�+o�5���&�$EZY������ ��?�oq�2v�l�˞�Z�r�,��&CFz�dn^�%yC�wN��/�/�dR1�M!Svk��\0-�L����<٨�+�@�;0j������^(�4�<�x�޶�MHĜ=��4��.�{ԍ���	��5Z���1��}8A�Z�e(�jv���d���������4wM�%�Р���4�{I��\����n#�b�r��~�������)b��mh�������m9�����2_�>Y�nyъK����`�؆�\��S-;����>ga���F�zM"��z�ٜ-�������B�2�l���풐����6z���pk0	��JJ�w�ai�_�/9�hD�mJ��ŷ��������<<�"�+�qn���!pq�����c"���72���YBfY��b k�b5?{R��_M
�:�(��N�B_穘/�FA#SLO��+��\�+��s�E�J"
�@~y�q���������<�#�i��7?<�ᒏ�q����V�ݮp�����}������u��[&Py7u�*B4i�)�b=]�N�3f+�@bt�Kk�m3�p����u*�o还��u�;�"�(��!�J�*�L�E^z_��ƍO_��υG�kn2�_�kr�y\pWڗ黾SV:�B{�D��IN�:`(-k��u�@I��><pE�Մ�$��uv6�� Fp�3`����G�O��gѪ���Xh9�w����_�#��$MO��r%�<�=�e[���r9Jh��0j0m?Va����=u�Ǎztۦc��'@z���c,w'�gѢm�3db%lF��]2�.�u-��N%�xp7��0��)�&=)�a�=���?������#� ��s ���B����|�d�>�
�V���4�lt,��j��\�wC�
�/�#�d2���7��X�r]���������ۅqzo�X�@M�LzfA~p�e/�+d
�;u�@��FȂ��R\�T�+���>�ǰ�z5)�(��ı�Oޚhmr*��K��z1�=[-��XK��y[p�ZGΚ����:��?�AC�1Õ �Ў*0�'4/�Z��T�wi�p��Lά(�=#�j$�'iz}RM%F�
�X�D^A�G�9��9�E-[�T�V;|��b�zW
�$���o��|�H9:�������	����8ѩ�r`ط��1���?��0�Za���sP��37菽9��"�]�vF4�IGt���'���j-��ϒ�U�	�Ƃ�<k�d�;����Ś�	��F���g��ko�+�L��^���V�wEv⧝,�`.H#Oقؾ��hN�d�3����hԁ��H��?n�����M�~M��o��!��N�q1 ����!I&ȥ�s3��K��Hd�oQ�/�\��-�����j�vZd���Sx��#h@�+�}	2`ǥ�x�z��Hz}^�.Haҕf�f�Aj�`��Y����o�<��vX����I1�^|F5��)��5L{�������羃q�43 ��p�0xjߜ*s�����HE�(0�N������;am����C@E�R, ��n�ҙ	�#����6� �⳾�c���E�.��G�Řu�L��%/k�+�q���1̇v���t��r���3�!^��?��x�K�cj��������~1�k���nd�R���O]:��-ĶT��WR+���R�2W�c}�ؔ���=���hO�C��A��f�k-���i��w6 ��Or��y���\9��6=+�n�i�\gݡ��|�7ŘyR�i���U�j2��2��$Y�#vQ�V�0��>�U�ԥ˯���U��bm�	�i�m=CӐ1o4���]'e�Q� 7���dEK��MT�z��g�����޼�>�:�pj�>#zy%)�������z!.չ���G6�`+댎�p!}�2�h�)3�F��U�Ow�T�^!����B��%VpT*���=��7�^�t�	*a�-���d��*�OV| ��=�a�y��9�.[$/?�/�������j�;�iV��(K|���t����@=D�W�a�^�|�����6rz���h�%�����O���	T�Y�ƉH����M���o*[��bAG�u���rK$��d�L���A�P�+�@��DF��t�ʷ|wՑ}�*` c�9�f���;���\����A/�"R�1:�(}�UF-�����(�o����'}��ѥ��ai!&̞5��O&#�s��\_y���n&~��ѓTi"Dd�;+�:�$A�s\���Em#]�N��r��������%���Τ�4��S;�(7��ɂ�{�F���8y�Ǫ_+x�ŁԄxW��H��ު����|Ev��F��L����c1z��7����k����J�w�2;{M<ի�Z�$8/+IR;�����lx����[���q{�Q-f�(CE���亀u���9��q�(z�F�&�#	3X��Iʱ�����<fЛ�6Yb�E��I��A+ ��֓GJ����n�E��������Kw`֪r]�#?P�����"B�G5���k� 4�m�\^��(gՑ*/�:���z�-��(�P�����d�6Ip�P\7|�=�M�]��ȝ��Ϯ��8ck��P�A��v�b�۹�($� a�ڣ���nY��c6
I��M�a�fm������O�ߊ�����Pɹ�XlxV64EB     a44     2c0��`.����� $0V��=��q�n�St5�`���7=ĵ�{y�;">����L��_g��7��"*��k*6�:*U�U�Q��5l�F��/[�[��c2o��ɯ;,���I����Y����o�Cjtn|�d�5��'���~�sH���V�M`�f!v��b��v[P�U�e�]٭�ف���P@E�O�E$�7Qre�z!�?��y�~�&�����UjP�{%v���=U;?7��&�����+;-�򧮱\�TpA Vnx��+�d��8{15�3����]�0V� �D� �>BbuV6�2���̿�2Ơ�&��r��ʾ��c���C��mG�\L_��a�d���������á����ȃ�&<��~�8�q��"�Mzt�5T��ԯ���1|�e��K����9��S�sL�y���qn2�zx��B8c^0oy��6����^Q+�[�-0(F^�PW��\K������eȏ��� B\<��d������ǖ�EU/��PSh�p�LT`C�lL��=���uDy�#@�m`F\{YĻ�D�bT��l�I����V5O=���&��v�U�Y����]3��۩u��&Y�VwƠRA�<2����!-@ڦA!�Y��c?;V��,6���ig�0d#�4[�UU1�],��R�Ҹ���'� SnF�I��h:P�`��
�R�