XlxV64EB    8c6e    1540�.� �?��y��A4;�*Ug�P}6Uk��>�u��D�c�[�֣�0�,�դ�c�@�{�I^�?��_����z;�Q����Ez��t��t��*��NLuOw���Β�3%'����'����-���~x�\��]�^�*�Y��3l��v�{��n["#��r�T5AFK��w��7ql��?}"���g�f�&����%Ә��*�0_�-f�*��(�%��u[�(Y=d�*x�?"Ϟv�:Q��M��=��,��f��G�葷�I��.����v�?;�!��Xz�M囅��p�x������w�x+x	D����E;E7QO�=���I�?O--p�V`.�aO�3`�|�f���{~gI���������o�<����z��/�]P���t�覡I�Z�Q�d��C���hC���b�7�X�YP�ML�/+�L}f��[@������ٙr���=���>�}��cTI��c�	��8��5Ԯ-�I˩��?�)9�B�j��&s���=u��1"�Z�R�'�2���^�=�,�W���H.�F������t�X�XףC$ˇ���W��VA����$ë�$��@����;28���1��D!*�S۹:
�;6����#�0Yg�TE�(
	_��H:�k*��L��
�������%�@�7ѕ���􈳻�\�6���8`o���YL{�ө��>5��\���f�L�/w+�>�xʱ��A�oO�q�9�v$�|�Y�MKwS�6*�6�NU[��̔g'&��f:����[�����3�� 
\�*t�(u�s��G� r�WF,�g��f�WR��vd-�l/Y��%ecAT�^��h��E��_z��[8���OrN�M����ҦHR��Հ�]��+V]��8��ʕ�ה-T^w%�~L�?��|'�w�35^̆�+p�"���_����|��ޏ5K2K�z>�	��T�Y�_��#A�H)�B��X�+�h��&��9	)�i!�J�U´͝m�'�L&8Yq��5nN4��WVQ�O&�H1���ns�Q��}%�(A�B�y�k���^a�êe��2F�FSN�j���8�q��	ց���fV	��7��g>��x�_${��^��7Z ���}kD�?a��:6Ȯ�lRM
c�-W����|�w�
e�}��?�5%OY"&�WH�8g0wXW�	=H`���{V�Q�ߠ�)��:\Z��e�:�+p	~
���0��h�J,������ɝ1�����-�A	l�n���f�:�XU4��}�7B.�����[����q��+jv6c)���ɮ5����#��n�GUNL�.H6�n*�,ɸm���]���&����k��R}(\�TZM\��~<g��t��iq�Y�b2Ħ��?�����'�C�h2(��hh��G��!v�?����(�>7(��l'¹���J��N�&���L]��+�x�O������(%!��������h֨�[[J�AǢ�ʽҚE��9��A�������E�;��IA���������!GF�|��Z�����G�X0���l�M�2�� 1L�e�uѭ\y�D�-������t�?�;icJg������e}y[�k��%H]�	�w�)v�i�Ur	�8/��l\��̀Q�U���j�,?�oo���)8V�oH��2��tO+.�S�uN�+�O�����-��2�nxD��k[�M�})�X����5�H��g��KDn���S}�3?�U�1��Z2�R>���[wWӒ4]����>&�Zpp��pV���%�$��s��5&�	�����B�S�����i���6<��r�ߣb|W(�sr�6%JE�+�̩��|������u��1}�YO�]���o
�����G�^��<Y=z���E���;�Zs���@ZŬ1��ԌA+/X�Ȅu-EN@ Cn��5z߃�q�뉔D������,5�K��'0BI_�@I�"����$�G�-�_�	�S�|�>���7��}��鲪�:@�*A.����T��W��г;��y�U�0�����#��p�2��۲�S����t�v-L�5���+8p��W�B��I)����o�r��Q-W�����p�i$��
�2��d��i�)"�Ǧ6���8����Υ�M�,��&�K%����ݜ�baDG��'��`;SP�ર�� E� ��ޖ���J�xZ���5�8������<l0&�kqU�S�z8���QT�s/~���`��L �����.��,�s��n�.�&�\��Ad'�8�t��*e�X�.*�����l8a�����?�X����cr�r��n�#�A��6���S.Np9����7(��/�s�Q`X�R	u]t�!��z��Ų�n�י��5cqph%��3Y�YV�őC�Cѻt��g�	�t�<����x��?]fwe7β�q��*���&8���_މ�q�RId�Ot
��G�C�O�uM���d$�W���t&��5�]�3b�9K~\�m�B��� (��Kv�#��_���ȍs>V{?�*=�ُ-[���@��"�'�|
CA׍ֈ¦{xUm���].�m�Ī�v»��i:���V��3� �#��&�)t��}�½N)oɃ��k/X���Z���J�xn/�޷���p�ߞ�6�_��H&a��&>�*�ۂZ{�Y�#c��B7����W6��:8+I��Q)�i}I4e2<Gm/�Ʌi��_�������i�r��P��~�h���*]2����L�'�)���x}��N��Ra����3ǕԷ�雎��,��xq��>�h*�4��Gē�<�.|�|��#Xϊ�r�4�,��0��h.���ڣ$^Ҫ������2j{l��@;H7LƏ�Fi�EK[�ϔ���ށ�-�I�ڛ������pV�a��is��.��&d��J�Z�樌I!��˸O��-v�%��2�=8�5��'�Cʧ�Z#K���FQ���`S8W����
�=��$�"���hu��fԤ����%��;z���ÿ��y~8��C�`�<,�h2�˴`��Y�6���3I㱲�v�=�_�6ȳ�&�ãb�c����B/�&\=��e�����Q)��+�����v�PO2᭶��pQ�����("ƞ0p�����6�
�2��GUyK�{cG�&�4���)�F���B�E�Q��`���~ɒٗPԹ �A����Q%��'}�F���Yk]�����ENu[��l�G��Nħ�����G���R�i3�|��W�TẏݴJ�����8�QK��L�p
T(��<2L�=��=�w���#=�E���k�/5���D܆,���TF���2$/�*Ik���~�����2��Cl�"�PV>���V��!�}w�bJ�
��K��N�G���F鄾^��Ys�	�����98���7w�u�er|W���K;H�'O�G�B2�J�g�d@LY��8X��w��N���p�G��<\T*:�ɐI����W�ʟo�]��KQq��]�@��)��O�o��ڗ�%H��q�X3nI����Uh�&�X\�ؾ�H �yI���N�V�Uj*F�����JFb%��,��M�Z�s�r5kg���SQ��\3)�!yf���0#,+��g]`T�c��� .Pk��vԀlf
æ8d��v�뭼*����7��pts��Y�/���2�d@����M,X���)��df�'���"�5"��]�
w ޏt��|ω/u���Yĵ��A+@ِ�c]�8��c�vgm�g&�@�,�k�7O�� �pĖ<9�H885��;���/Q��5@�e"B���#��~Ej�4̫�Z�':�($�5Ol�#	M�v�*s�1� Q�934V�)$E�� Z]1 ,r,�*�8Q��\�ܢE���ωl�n�v�"ѿt]��X����?��6�N�`rzϓ8�Y��|���������wh���?,��	�8��2R�=���#?��W�����R�t���j��x�,���$G.�j��)�9S>1:����	�f�J��Yf��8C�z	?-l��S���O;GlOA ���Ҷ�ڭ�8��vvG��󅣡��~�a���7�'=a�:fl����2������+� K��f������S-�����p>
&T%�Vd�OeY�5̨�̹��2�Jܱ�>G��2wg\�;�q��æ%q��u��tz���AC���'��=c�^KP��?���`��xK����Z�z����t���s�v_����g LDh��������g[�����_���: �5�E=A����g��Y�o�i)��;�ӿ�!��,N �FE�ݓ���M?s����;O�� ���E��������z����el]MR�h�}����p�+@�J2T 9V�s]�J�'�Bדk�k�.����g��6����2U@���\�#}m`"D#�α���7���ڜ�@U�9�y�&S���䂅���r���W �4�v��O��ʄ�S��-��$R}��I�i,��E����38��=�|�CH�wQ���^ֵ?j���MD�w(�W�9 �$~j�<˻���)�J�[d���\��͍&�~"?��j��p�z9dլh���=�ę�gy�?jcRn��Q��ۜ�z�^��ۅ��۶�gSxƂ�!$P�)�5��H1��p�.} <+��������2�	l�͈V�t�r�uz�'�������cd���5��x���Y�7�y�����\Lط�ڂ���r�*�)e3G
�v���aXto�SP,;�S�lfjj�lE�_��^e_a���㝖�"���Фp��.��1�9K^��K�;b�А�S;�;D~R߃�ϗ��لk�s��Y?���F`�P�yGb�J�7�v(I��BD����x��nN{�:�[E�R �V�D�����z�_�mn/��^l]R�.�pͦ�z��!W�X҈���qup�!o�&=q�b$�ZȵZ�S)K>$�$}����b�GA!),!pP��m���bJ����:KK���Օ~W�;�Y���/j�4�RC:�]͕>�0@��%͕	�QU��>劮<σ+1���F�y6H�iYF�_�%�[��h4[%���z!�Mn��o��7vJo����9��{��Ċ��Uܵ�=H0r4�K�8c9�\oL��T��Q��Q�$xh;U���B�$��<�N��U����u�N�~9�Gp�z��}�Q";5�׬q�pW�O�,�f�[�^�ؿ�	8^���Im:+�,���4T2F ����ߓZ���nd�w1/�t�k�x#3��Ft�A��`��$���Aqx}��d�+4������by��j��
P��^4PJ�&1E�Vu�B�z�v��;gЮ���	>	�pt!�<X!c