XlxV64EB    4110     dd0v�6�
�6��B~7���[`�.z������ �ylp>d��v��Fݳ�<�j�_�ХL��n�8fu�ך@��ʐ� �Q)S(|R\H�+��O�d���@����d}���>u�wܬ�
�`��D���w�9���X��2����L� �cM�l�`O�6'q,��{��� ���E�V�ѤF3g�A���e0�'�ڸ�N8�MD�s�����̤�:|�+dm�g�V�D8�p�7"����4$ �0���c����f���g�C��$Z�q������9�תSA�9��>d,М1w�&�@���R����ٲ����� ԑ�����/������|�g��M�ؕک� 4�җP�?RfL������>o�/"}�}D���#�8�Q�������p�J1/����-4>�'f�
�N�![CD�Βr�\����s�� 7���A\3)C߾%�%a0���N����_S���I	9zëj� c��8��>�|�w6���ؚ�@i��gO*z~&+�Ga�ǲ��wܭ~_��̥��n�S���r������N׍�z\���m�J����M��ׅ`�"d7�
Y��&`<¸����T�ou'k���vY�m��ШV��}�L��|�E�DE���":�b�,��ޤ�9��
^9��j��s��'����Пs�O�`�.m���Q�'k�s�d�lW$�:%����>��(�>����̛�#� �?���?
U�A����(�ɧ�R{�2>��ʅ������o��d)Ȃs��j����4��&���n���Z���3��$�DJ�-�ۊ1�w�m:�;@��j���1��nV�kW�!Q�]9���Y���馻��7��/D�xC����[.�km���d��Lm�+P��̿w�c���Tt�wa"���V�0�
;Ød0`��TB�xLc�Q	(	�܂��h����:�E�Ln�/�ks0���_'�='g{��Vz8��~ǧ��m륈vĄ��I� :*b������;j�(ٹ���P#'��Z����?�����8�*�!�� �3mu�2��r�fw:�+�����KT=�8lx����D|���Ɣ�+�w��}��X%HR�{تg�&��t��|e��37R�M�SN���Eʲy�=�֥���ʦ.����&+����������D��&��'�@jg��"�:R,+�K}��c�Q��T�~��'�O�i���3yp��-V"LJrX��-����P��M'���1��Ե���j�s��3S���!�W�������#���#=9�U�I�b/-0ǎ��`���^ ^X�B Lx��&�t&�DqҬ'��5�JF��-�
���Ǳ{뜇��ß1pY�,D���6�Ѧ-g�Uc�1�~,xpw��;a�v�TB���F�
q�0ܿC��Ͻ�g�\��ê��Ӷ�y���U�\��}��祥w��䰡�E��Znځp?�X�1�W>E��Im�M�X�^�Ƕ�XjRr�P�E9��jۢ���)0�T�=�~�ҶB�#�*AI�
��F*W6�w�S.h�W<�|qh	�}a���8����(��z�`y�2srp�xj�$�}�lm����\]P$���U����f���#��`썔Vn����E5�ZPt�v���K�LZ�`6�ו����y\�a��w��\x	���Z���:4�#�A�����zMG\����F���K�Q�W�� �����q3?A	ϊ8�%��v1��좟�����C[��=�DK�>r�����z#y1�	�r���l_)O�H���Hb蘳�_C&E����H	c8�N�|�녋�nY~^=�~D������&@M�y����]O޴��dP��_��l���,�~f�_�)C$ᦳ��fa�@a��7���{�F4qh6�=��w�8I�nI���ckZ��S
{��yfY�4�q:�j�]b����p��s���'廮��yP�J`]��V�{}V�R	����U��,�d��6��)+(+�Vc����P+[)�2e$/՛ZU���<�|17p
��haa�f�-���cڲ6�T<|�^����^U���ڵ�}<OZ6��,e����`	G���<%l�*뺥�0�,�dJt�����n��5Oc���AЍ=�~����,=-��\�~����Z��a*��:uZ�0t]�8�^J��6�*���=O��U#gz�v���Q4�Sqٸ�I�s�}(7�
���
hC������p��;�ն�B#4�z+P��������Qԇ�(g��UH\Վ��&�Q�>�8cꢧ�i�Vנ��~�<�^������l&� ���Auq&��Ҝ��r��\ڱ�<���x<4�$�x�a�"=S&��:�Z�@�1>B�M�O*"��ܶ>���2�蒿�+w�K�e�2�(IL#�;X~Ȧ@��e��˰k2?&���Ƴ�#���C��<j�D"����2}��c	�,�t��/{�j[B?�[ǱhP���Jnȷ��Z���Ĉ݇ʵ�6��"KL�!ÎT����u�xj=m��$@�߫����X���\$��Դ/�S������zy-b�,'������Z�j��p���bk�z�Ǖ>)�u�Q�*�!bJ�:��J?G���0�l��m�64rf�������2�Y���1����7�QZ,W�٘n�榏�'�vB�.�H�7_ɭ/���ѾAL*@��=:�?OZ���,��|bАr|�'���n��q_Ģ�3�>CO�hl�#�(寵�-K���&�fտ$x񍥊�����V���;�ϏT�y;�'t���X��.��r���c��9�3Ha�Э������@���*�B��*�>MU�Ն6ܸ���Ȃ櫯��)�&�Y2Q�f�Q��W/����
�G��SY���>rE_Ed��آs��7�0�������E�1�1�%��ހ淮�f(A����I��)���*���{#�p�����Z��^�K��0:���cЮ	����� ���ȎE��oB�_{N����X�Ñ(Qh�S�
��}��ޝ��j�5^��WeRN����lY�`��3#���XD��#���g����o���Qv_�A�f�w�}:�h�x����i~ˣ7���M�g�u{�P=,x���e���+�ly���T�*��C�
S�{s-�s/9Q��Q�iik�m]��B�/�* �B�A�� wv�+4D5\��g�쬭x.QDb��Q� ���C�4L��pXׂý�I�6��I-H�������x�x��^�֏����u���-D5$�P=Ψ��W͓�H����"e����E[\N V1�Ҭ(@Q�G��nE�aVv��i�R�8&����e���f*n�׈$�:e �h��q�TAy��ƶ�U?��:s,C�+/�Ā����vEÖ�l�Y]Q^�����T��gI��B����N�_D"�^O9����YT�o�k���[5���)���t���|�o��7CC[�]