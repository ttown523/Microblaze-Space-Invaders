XlxV64EB    1f15     a50a�ŸV����eoy��vA��O-Dd/����!�Fx���qIv��K6�����[�"7��h^��/��"�y���IV�yeK{ƾ���~�̍�������J�,Y�y�B̥�G�sR���^�7Y�":�2��w��ÓGSO�ȹ���X(e�!|�ZX�� ���m��P�� �`�����o���l?σ�>��@2��)��@����	BÃ�Ԃ�ʺ�3]���,�� IPзN�Bg�ud�&~"�b{�3�o���$#���-�T"�������R�y�����ۗ �m���H���V�� �K���L]��OV�������;��8 ���Tț�U?jM��s�������=�|�ݘQ˘7|�7!FƯ��{h��8����u�̻b�- ���F�M��=vG����}�V��B��2�&�"<�� �֌�ω�,fͿdіK^�8�R!4ƺ����l�[?��ۧ�=�ẋ��׬��#A�W�u?c�/��(�$3�����Y��e�L�E&B�`��µ$Ry�4X8s���E)j*T�b��y>����h| �������k���N�����a�C}X����N�
� ���1��|H�kH�n��?P�p�4
st&fظQi{dW���c'��	�CW�Т���T�Ca�kj\���]�M�����){�"]Mc� <����T|�D3�@�m�j�򲺑�J:W�x�H�������E�
��[H���������~�>���b��ۓ�O2Dl�c�҅�
�W��R�-�}Q��xS��o�~�?CRr�E7�y��Q)_x�8�a�<ܟ�)�I�K�e,Dɮ"A~���A��]���L�d��or��{bYꈺ��b�+����������R�ǿ��C0�}�'�H��h��o4-q�U%�4� ?�|(?��B�߃�_L���Uft&q��({7i$��k���:P�Ac[�P_������7�7��j6l[�K#p���4@:��zʑy3����&.&!��ʶ<��q��C̎5�TP�ѲW���rw�TH��B�蔾�o$�<�<�S1e\���r�V�������DYMw�h��#�~��x�������L�I��g�>�-�k�/�_,ޢPH	IjpA|��a���'>Y8�.Y�HWB��xDJ��Mc��A_Wqz����ڬ���U+�]&�&h@���kG2o�cbM6�R���u|� N�y1jM`к�<��G��ʙ�2�u�~���F�>�Ո�vb0�����PN�i�H)����d��w<[��-�׌9[$P��p��&Ȗ�z�ՆY�n����[�|%L^H��	BwF�l���R����Ɲ�C�w���ճu&���r���6���������9c��Y��N�����S�w���7�
�R�f�v�����P1j5@Gc~�ܵ{�K 2U��+�$w�da(V�$PL�<��axe����hd����X��8�c�d�m����ʏm�!��'�8$�����ׯFo�Κ�����@ւa'h!H�Ϫ+/&�����bS�S^�,6�(�~�K�1�H39o�K6���Ap��e�-���U�վ-jC���iY�.��]����u�R-S�
C� υI:舱������Y�d�yﴊ8����aHr������R���V*�P��z��BW3�G:�����yyD!|�^��.�³��=�o�K���N6juNֆ3��_��vAET��-�fz�
��J	�g�1\�ڒ=����m$��;�s����P�LV����fq��\�#�z����х�Wy
��`���l1}�N4:�J��$1�	n �E���l.��t�<��� '2wT����o�fKFk]/僯 ɡZ��p�m�Ĺ����&�������y��{��U^}RU �%�e�}K���#�L6b��ԹG+���KD�h��c3�ŭaZJ	�U⿹֝wYb~�c���.-o9�����f�=���Ý�J��Vu��.j<���d�8 L޲ ��y��u� ��G�U����v��o�wײ);0�?K�2k,܎)��|��꾞��������s9g��m��'��s<���	 ��&��US��o(�=��y���e���H�/_4Er�~��L����i�MC!@Xm�(z��,\8�ŏ?�sX�g���n�'O��?L�S�?O��z�+��xp}w�>�*�+X/�eg	���$�ή�fq:L�e#S�Q&�f�G�1�q-9�y�f�ʏ7�f�4�cm�<��ٱ<�Z�9�v�3O,���iS�P��s=&ұ�XOEG���B��{���6���$���^vf��	�
�Q֤k�@�?����6j�X��2HR;��-8N��u좧�-A�m���s=Ů�9m�b[d�G�w�r���uS�S��&��;�]oW��7�5�u�f�b��
Ci�OJ�@ʯQjB̟���l��ȴ��INm�?�l��80R�k�� K�G9�	C�+��>���ۧ|`á���S�M��3�`۸W�Lo���$����HcO�������`��0���M�x��f�G�_��W��Yùvl���Ϣ����"