XlxV64EB    168b     8b0�q��ed�˺��
�WY�.Zs���\|���K�_����Ը"��H��ŕ�`Q�h�,'�v_Zk��z� ,���%Z9�Y�U�t��`�ەb�R����̣������4l�ݛi,��dB��(c>���0gy�e��TPⵚ�H��`0r!U=�<��j��N��Q��sx���������;ȁY�M�.�Ҙ��,[y%�;"؀13���G���[})�N�a�,��赽����حDŎ:��⪌� �����I���sBadu�ShCT}�k��U�|Y�l�-�s-�ߘj�+S��Ѳ���g~rzh�����MHVg�D�1�?����3d�qR�z;R�;f<�W|��L����w�g<7��f�5�����"���ܸ�,�	@]ߢ�w
��H�d�\����[�9��럢��h)�Vz�I͛���P�h�-	YO�x�h0��ZsL��}
�#�rP#���`�����	��/�X��j���V8�Y4��G�R�^�4?fŹk˒4��{�"�<�����UR7�x�.h�k�C��CUaA�'^)m׆��C�^�A��I����	�w�M�e��@��E��V�+���uT:�Z���I%]�焔�᳒���d/�j^��-��]� ����{��K��V���e	[��b�&��[�P�@N�ED..W�s��F��0+Hw�p��I]���ڪ7v���2.�	ҍ���ֲҴ�&{Q�c�ILYaQ�)�m�rM����0��L�1r����v���H�_:�;�H�5�x�7�OȖQ�Ki2�;���n�����u�<,����ż�D��K5��0��Jޭ�h斘ݸ�^��G{�$;?[g�#�j>5�2�=V|.��=�'�,��ڙ����q���~Μ��;.o(�&��(#�
�Qc�Q�ҧ.�ׅЎtCM��0��xU���½Z��Q��w��VN��TkSB��3�㪡��?h�X�"�n��t�!gUv�Ѥ{��[`��)�(�hq�����X��^�RS��/�7�]��s�B/AF��.,u��*��Фe�L��x��d��� (#df�EޔO9�J�۴t\����fpIJT�v�[���<�*LڡP�o�o�e:�P��KtS%���z)�|�@�~G���2�w�u�����Vn�b"��Ma�k�65�)�ۆ{v��p������qk���h��Mң7%d�;��V�\H\[�w+�b��C���1�m���Zg}(p=��9�<v��L�v�':��	�Ӽ ^���� "�X�ᢥ�q"h���ƭ��W�5���_T&,��vw�o�_����K~)�&i�b�6}f�l���H�#8ۚ ����.U�$6�t�)��^�j�"8�'��^�U�V�2�c��-�y��9zT\�=h���<���@��h �k�B�2�g<�ȧq�= ��s(��8(�xq`���"���oK����%��*$�\�&�3;.
o_��U�#���ŋr�*�T%P�|���Nq|�L�r[��㭳�7��4s�v_�L/~n��m�O&C����,���K��Ù̞aZ���mL�m�z5��������k��B��UZ0㥺�¾���L�����B�m7%ȒyX�Q]�̦�X�#*��FNi���H�8dLIb.�������0j��]�����k+�Ӿ1���`����"_������½���4F+��u�\�VY?��H_B����{+mh��c(�?�����6�D~��^z�\vIp��AJ �M�B2l�A������2��
+����3{[-�H�px�۟d7?�|c �����Ү'���4�����{Z���ı�����������{�.�ւ���xS:�8#�Z<7$N�@�%(�#�n<��.i"V����B����Bj1��:�������}}o��`��M��tzV�^�����W�������v�,���4a�6�օ�\��A.Eq�h��<��G 0�����}`�>�a����M�1,5 iXc1.2�KZ/���,djF&I7���5���K�_"L��jxܾDk��yRb���j)o� �V_�����������{O��S�W>6Vw';?+c_�T�����>�2^(�xťF̗� �M<s�N&O�Y�z�(�Xtx�w��7ka�0i(���)B���@���r����&��$[&���MB�������-5�կ��n���S