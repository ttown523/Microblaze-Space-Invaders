XlxV64EB    c9d8    1a502���:�*�\�W	�p������1�����U$���������S�E]yKji�A�\7fu|[�g1�u��ji�\��0�2�߄���T"ʙ���p��K�N��	h����k����z��`V�i^V�2�>D �9{�/�N�PVmˮ����<D�[%*_,g�䢩
r��l�bq6�H�E�Y]�oA�#�ѹk�h�n�q���cv��i� N� rX��*�836���~@��	���W"���(>��36Nz�w���'�9����{�I;v¨�'NzAk{���YL��*�	�Ŭ^x;�����I�;�c�<������ّ�id$m�^�g��nգP�=��~@���[)��?�����"����|�?�x��X�
���KE���1=�CCC�I��L��-���T����"��� �J`8&��a��Ec�(_h��$�'��:D6�� �Lb�r�0q,����;�qn?��ۦ	���� g
�'�[r΅�]�����os �	�����60(��L"k_Z�}/<�P���+�X�cV�L���E����ج��J
	<9 zb��ԣ�'�ah)v�������f?B�by��tO�N�(����8w(�`��5/��f�p}#�,�2�C]�C�c�G<ݮ�����e�Ia�n�PxM�q���x`��%,���A����9ֹނ��KB�qR�C���,��YD��cDҋ�E��Y��C�Yg����9^Lt�R��Q 3�'8�R��s�ƺJ���F��V�\��o\_ȹCH��>	w�yO�ᘻ�8���^{�¼eW�s����M�ɼ&+��E���s��g�f�۫��L<��!
3w�2����m�T R�4�}��%7��d.ؿ��ر�^:�论��rH���]�X����ڔ�X�������"eX� ��G"��֏���E��Tp��Ѷ8ܱ��;�K��.�
��,�܃h
C��3��a9F#i��萅6ڣ�OBID;yl���E����q��^�$~*mc"~�.f."�tfF�j�e���
^= #f.����d��B��Z3��)�y��Vk~���fplt�*Ҩ��*�`yi�L�nI�`?ӢT-�Yל����3%ށ��
�<��0m,p� ��Ρbu�"霮�v�*h������^�F�<4LmL��X=�z���ߟIX?���*�'_}�"�qS�8�d����i6���<w��8�����s@@y?�_�
�&D9ړ�`��(a�r�e��׻%�d9ǽZk��z���%��Q�M�UÞ�� �"�����>�ȃ��"}�EQ�n�	��q���P*�jd0�I!�R"8�80b A�0��������:x�"����I�}>.K�k��Z�R�O��F����l(6�%�Ҝ�D8����(���"=u������e\q��2��;Fk�)�$
`lu����:��yC!�\N���H6�źĤC�c��f ��/�SN�����V~�L���&{2 ��k��ohI��Vc�ݠᖏ���pq�
��f��^�a���^�֖��K���b�JJ��>���S6���6ĒI�o <k?�'�$���3�k����iN����'����ˣ��/��6��թ[j��J��+
"rX/��D�΍R�P����T����z�\��j�E``��Y2����*�X���F��c	z����iĂև�j<�<�dA;>ʼ��W3;Ǌ��\跺-�~��� ���q<���l�1���u�[����`�c�y^ �M%����"�/�������	ݬ���$����v�n�����G8�̋$��[j[��/0͉���_���g�а��e	ޜ�@?\����P�P��'���=���[!hլ�s_���(�Or�s}�Y,��`9S)r�zg�]�(m�ck��Vf�Bc
/ʰ��_VӉ���%����l\AVe<��L&ɽ)�#dX�h8�C�-X���I��;7��2��ZB�)��r�l�������d���-� ���?��_Y#�^O��έ�J��kKX��.���U�������+j\��]�żR-ɉ0�pP��!�H:��7��lʟ"i����`=�f���.�Uv޼Z�<�|�_�i7A+cNY����4G�a��ҙ-<���~:V����^�hU�w�5����42�������~��X�`�x(��fȿ�?n�ŏ�E��mK��?���c�[	7�`(����
-*�Y��[�e��b=rmxK���l¬�� 2��"J[	���6��`��q��c� MM#�d����	F�=��*W=q�d͝���%n�aȵ�6��X�TT�sz�Dި1P�/�U�Qr�H�vl�K�g��ɍ���N�R���m˘�h�2�Ka��E�z���K�	���Ix�E������QA��D{3Q���D�+�Y��=y֫�l�Z[���Z��*?	��Jʋ�2���@����4cs�YyY��]�������<Iq�{<�jy�8#��~
3��V4k��&3Hޞ���:B©jR�zuv�=��#�D#�m7d���S��u6���݌�qj�R>��|I�͐,��ێy��0nZ�/�c�g	Թ�a�
�/�.��a׳Y��F������?$�"�Xs��´��^N��� "I�P
���Y<����3��?cPPLUJI�G��Yb�팬RN [��}U��}?�V�-[ ���9l�
��ם]���h7��c��Iz��'�ne\�:�����3A��G:KWF΃�6�WV+BQ*i2<����[����������/��=6��3����p�.�	 q���@Pq��w8��)�3�R�&��-�0���~𠗈�P {"�¬g���_ݿ��QN
4�#�]���.nb�L�I���Gh"����	�z��{��<1����ᢙ�_	,E�˒�$Ŭ�ˉ��0��u�����)1'I��0� N�0��e���%��
�:����#��F�)kֵ��T]�D�����KN" rs*�ZK�.�0[z�'kqɟvy����$9G��9�x )G��H�K�'?�оO��o[_�n�طN2�|bR"�,D4���$g���եbɫa�=�[��7b}xc�%��|�[��*$^�$wKbg��n�N�:�"�����fc,��"GW������;��]�A�FWPeW����P0�{�&��>*�LoI!�&��\Bh�x7��..����K��h��P+��GF�h��9�al�ّ�¢�_e�*�H���$�? ���o��h�Ŷic�9�w��`��K��+��w�/�`'�d��̺$#r���2�^��%C[Z	�g�<|/J�Z�������Tט�3�՚�P�	I_�r/B��@��#C�6o�r`sB���uRk�B�&����8dF����Mtki-�z7�F.��o��9�@E���\n`P4�Sl[�Ee�\�8���.��K�� ֗5ig0�"wI�Q���{������4�<�°���[E�)����0y$Bs�r�&:����5��t�ΌF捾�=#RAĭ.?��rC�����x�5�A蝩;�rU+����6;�
e��A���G��H�b��z����(�ψA
�"#N�) ~"$�r�4�C,�'�TYvة(�1��O��[�����;�"�VC��qr�G����9��+\��pW!�_�tHD�`���K	h=ր[0��]���p��mG`�:��H��=}�j`�^� �WW ����Iꟙ9r>D����4R��T��>b�n<��Đx�HI��öKy���R�zm(9{�@�S�9��U� $q��)!\#����-HK Fux���v
�m�$����J��o�y����W�ic� Ȳ�u�%tA4s�z�յL]j��,�� ��bw�>��R��@���pn#[A�3�՜���)?Af?�_����.+5�]��D��<'KOcd�ZR �Ch6<�J�ο���A1x(��P{LP����g�Q�t%~A���!���W%̆+c�`����iȬ�INeǨ,��ng8|.jZ�-��u`�.�x��u��}��ت�������[��sy�/�hAÝ0
��?&"ح�D����7���}��������hrC'�i�L��P��z���ᅪ5U�??&��ϯ���*���jG ^�tW~����5�Xx���"�����׀э�7�W��6�.��駜�2��s��#�;:���I����K��`�h�ř,���12�������ӈ^���oӽ���f�������V�[���� ���i��3�x�KFɼ�4�<{�QXrkW�X�JUc� ̲1ċ�_�%0=�%�l�,T=%&���";�j�C߲2�LP�oީ��ѥ?G����$�1�_��6;[��M�m>F 6���s�. o���زS��D��f�iD3�(fpͩr����h�5m};<dyau-5��8l������[�2i}�4'$��~|wu��a���� ��z0���$�ݤʲ�v5���{���?�*���X�e��T�e�M'7�Jm��;��"�K(~�# �ur��f5hELe��1v��9b-�ֆ��a��1��B�5���h���Y�p_M�Yy��e��^c1�|�L�N`�A���h� |��\�^�����a�,���?�z�0+Jz��.s���	�S��wxȀQ��b�hV�@v%��>|�BOϒ��A:�<+HH�a@KO����S_�!	H$\�n^�u�����/\#�SO<�8ў��F .����⩹�s�nyRT�^���J6�2�7>F�O��W)�a��\���[���s�<~���N��ލf�S�
j�[�ȣ�����/<S����n��B��ˈ�7@�"W�a ԧ~}
!�Bɬe�5Α,��^�*���_���r�V�s|ݶ2���8��=�9�Q2�m�ޤ�=O��@���/+o:P%hs��y�v�o��
QD�e���$R�&�|�8��o���j�`ꐖ��D�W3���w�u�vk��@v?���3�~ ���|�^}R���H�p���	^\m��Y��i��$؆b�d��{
�a���ZrB��R�7�)2T�� <D�3�z�R�?��DT^����X=�w�)�
��C��	l�٧�<� _����Q�\�� |�\�|x��}xSv�Z_
K�9��,����b`��sF��bq�C�K�H7z+��-�Ѷ��G�XG�f�����3���Cky)N?Y��{��i;�Yk�?�?��?蕷"��M������3ˬ���M����^��X����"9��Xߘ�HmM��6�:/(�A��E����et�����\0����l���(@H؀Ău֤g��m�<g�E��ӂۯU�T��.�o�v��)�i���M�zL-| ��1�:7��%ܒO.�'�L=�1΢�7���v�T�����WCmy4Wߕ"�����������R�3M�'M]�|�'����1�����L&�K��1j*z��d��{"
Jߒdrd�tm
{i�K� =J�� dLr�?1�h�B�;/�qF�� cƺ��2.�E,#W��m���m�'��� <Kv�T�Ŭ�~%�WڻXU��˖�&�� ]B��'G���K�/e�5��q���U[O�U��8���[�����U��#l;k����\=���\d�lI�x6!��aݑ���U��x�|3��(l���|4#����s//�)b_V/�K��� /�9������~��$�{]�&�Q�eſ�P�bGE��L �L�z*3q�M����;k����
4����}��D�؝���=N�M!��A�����9qɻ�8���.��4� ��\z!A�]��B|;`}�x�������~��	?ώ�f�	1���!���A.��ײu���|�\�?4���NSEV�⴫�`���zC��ضj���԰�"�\΀Ç���/�W�非���%P��E�]zP59���~�l͈��:�n�3���e�L�SC9����w�Y"�&�k����/���΀�e�qKgg�_��64���;���ټ�<N�e���56킜��%D�y���~�W���G�q���J�$�t̄�"�(����e���l���W���'0�@4���
��,�<�7_�5�� �S�Y8�h���v*5*_Y	u>30�_H֐P��]?J(5-�L��9����đ��}�����\�.Q���7��Y�A����Ї�޽99:K��:�X�����6�U�:��� �<�ƈEa�Eg��b%�_�9���КE�ކ(m���Q&�}	�:�~�}�"8����U��'+�N�]\�be�*�����+�.�Û�&V_���~��BDY&�\�V����jw��jq�׍]���cܕؔ�a�S��-�xLU��7��4�xKR%},@����4Um*����#�W��MM�l�3�ܥ7�����ˇ^�!�����Os���
¾�_F� |�Y�#�&�N�rMc.t}�ȑ�~�	De,	��ˊe
���%,"O�gF�կ���0�⺗#�&�/@KR$؀@c�L��O�M�<�1��F��_�E�2��X�/f<ԩ�u!��a���Zs؃�c�H	l�:�