XlxV64EB    1feb     ae03C5�?�����2��Ct�h��/�\oU���G2�_j�N�Y�$ $j�gE�r+��r���\s�m����cqD9�v����b����vh������<�A���@�;�*��re�!�\��������Z�R��^WUB�8y�O��50�f7�#[�μ4�~��R��	щp+;������'Au�&���N�b��G�xM����u�j��r�X�5縭\�X�a���Y�[&���,���)'�G������ΐثY6w�+����e2&�C����h1"��Y{l���j�@<B�!�N��W{� Ѫy�� ����1'K�]Uآ��WI$LS�c鈩K��_
.1�%ɕ����3>h{f�,ݞ}їZ���:��<��J�������6<fʴ	�u׍�v|Z��gŉ4E*�q���NjI��
B���ؤ<�C�r�a0�cwp���ч�]�q���
�$���Pӎ�)�B�}��Z�9�e�6�b��ɀ@�
u5�k�������%�d �NU269ŗά�v�Pl�:\�	|�
̳:�Kd��#?�z��g��	$��uݱ }�<�QC |� 4��Z��u�>��E�C'���]I�.0!꾳wkG������ꆣ�*�W��ݿ����Y1A��V;=�p�.K�Qj�]`O�Qq���ыQe�|��\$T�$���&���1ۿ�YSr�Ĵ�5p�!�ݓ�ONkM�`F7�Y#��)� �g��:�M��U�rkx�B�M��C����B�әKf�a��9D����:j��>������n��0���%�8�w)��*�hg�Hӏ�Y8r u����;I͟aYPNΔ�F����/P���҉ݑ�U�/�����ۉcׅë)"î���<�V:Gy�"J���a��}�1L\�K2��V�	2U>	��U�+��}�|a�Ěͯk��	���lOa�_���A��Q���% pLF߁��t(cx:�Jߒl�"���/7$��[Q9�_�����ٮ���s�#����-�s���P����&+%;Y@#`o-��8MŎ�3�eQ���a�-,=�mK���>` 0V�׺��dp'-)F�����cA+�; �@���iR��峞�5��
�#�P$p�š&`QҘ�=5e�kQ���OM�)�~�lYl�6^�a��Gv��-��~���K��%�i�q)|Ya����vu�Z��2	�b4=-s<fe����	[+I�����,�*e���c����������6^Q!��Ň���Ydj���0tUm������ ]@q�<1L�i�[R4}��ӭ~8�b/�a#���JLrZH`_;�mdƗ��|t��2����4���cĤ!*�n�Cm2~ �"�G��8H5�L-��n78I�����<���sEY�.χ��R�Ps���y�o�؜�]{9l��������jAͧBÕWL%D_λ�Sʈ��k$	&�����X����n����K�e�p.l�%&��ړ_a�H�!֚l�"��Z�NH�,��L
���W���6ٙ���;}�����
!luB��~�8�����ސ�5t�^���v��x��PڲzA�޷,����E�	Ek��앐U"�B�V٣��D̻^J�f�'�T���P�j���l��o����h#��h����U�=�p��4%^�ըVy�(mju�<�D[r��Fm1]���6vg1�Ff�i�ᕿ�1��-���+�(�x�(�N%�æA��y|�������c8fk��dq��J�(�Ѭ�����5q��mN��7Tz,mΐӊ���gnew��)�"�Tm@|��!v�π\O?Q�Ƭ��"Y��T��3���j�K�~����;�(��Om
j͹gb� ��Pڙ&i�B�QmA���ǖ�.���G�! ��7X��x�
��(P��W�v����r���cf%%�3�0��o��	�
������5^�1�A���:.'�>dGA}�ټ�wb&Hl���횺�[*E�a��	M�jJ�Od2�Q����a�����K����ֹd�j�⩦ʇ�]u�32T'W!�)���#:ު�b���ã��ܤ����v:p|��=����\����QU�3h�,�w��ӕƞbd��J(t��a��8G���͘F�x��cO3�����!�l���}VWe�vLChpQ��K)=�A��$[�K��(@�^�;1�]}�xoU��:��C�D[��K܅�#��5vh�Z99�r�1$jѯ{�;m����a(���nG�k����W�ߴ�
7��'�+�,��k8��s~��{��Cjy��Z�?�a����3 0��D����Ժ��T�~�?�vuB�,�D����~>��FP������&A*-���M����y�uFQi��e��a7M�V�Ur09WC-κ <n�5�;U���հʢ�ԦDg"��'P�V^~� Z�)����	__.S��QIr���S˽�}!�k%B�L��Zς��\y���r�0`�e-W�]�Z!S?���I��r]�A�ߔ�9
R�<�L�429��m��˱)���r�>R��}��t�c���O�R�@��QϜr�c���m��V��d�M�R�|l
&_�>#G �Od����q�l��0��oX=f��d��� 7aϾ~���P�W�y�z	��0�Mo�Qr�'i�y�����m(hZs�|���-`��}J���	��pS`C�M}�3��+��