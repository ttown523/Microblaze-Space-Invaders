XlxV64EB    53e7    1140%�g:���F��0�Q�F䑧+���}�*+ay��Ӣ�����}��B
��@.2j�,�E�5�b4�84җ4Ѱk���b�;`�Ы�	���\�rr�Ŧ�H�<.���p&0�x��U<�e� �<zl�Ñ�A?����Ol�h/�Z��	�2��q-Ñ���o��S��s7�P�42S��O68<��ds��W�8�f˹�#����ٶ�~1?x��݈Ws��n���B�q�p�=݇}%���A�!uZ[��3mG�.��Hn�hP�9սL]�g%�Q���*z�hU�GW	�<X��D}��tA����9� +'�,0y��|��^��fZLI]`9á8�zi���V���`�I?�ćetM���8������myE�8��v�H�{����Los\�Ȳ����hߨ��<�1�����>7gj$zh��;�k��@��U�J�����s�V���:"�-���=���W[(�x<��5'a^ ݙܸ/��W~�c���_�Mi�%�v�i��0��I��8��/����y2�CE�"1/N��s���.�A��7�� ���Q�V8se�#��b��'�F$H
y���s���_vGQ_o���o�_&�N�D�`����K1n��=��7���˳������zX�Gf1ȵ���52���$�<�Y;������--so^�#W!mˬ�jz#��0���|E�8�K�\���[G� 6
W&X=TK�}U�D)d�f��_��e��𓕝R�`;�0ա�1?��1���Vqs��3���ɣ��ϫ�B�dR�k�*9;��A3�?�vH��$"��˅y<`��$^��*�@��u!�kId�,D,��G0��������i0W9�����^���y�Ш�sb"����^�&2+����:g@rw��7maw =L�Fx��tLq�Z�6Eo�o	�8N�23�3"�`!�W<��}p�e0�s汾�� ���:K���k�0$B�� �YT����^}(%�Pѱ��XX��>��l7���]�w�/�MK5�L		IcE^�7���*��c��q,ҙ�/��s���%u�=�z�X&�	�__�ׂqQf;���1�d��0!�W�w�	���$2U����_�"Xى���̔o[,��p�u-}���BJ�>y\Ji���ef�(�[V�˞3�{��ŕ��8r��o%#�H�G�)G|.��k��ckK����y&/�� ��V�f5y�2�])�f�Xp��䞠�����"ط�i@����)�����ُP���Ujf���&Z ��R��߬�+�1ɹ�lרFmh�XM_�vCJl#��m�5��Tl����a��-{_F
�V,�/Z莇�}��&�D��ݬ�n�$ɽ���"z��2`pb9�E�1+�=�D��2����30?j�~�D�7"�����bm�9��CF
ET��Yd{Ǐr>p�5�4�h���.�h�B�Af"������ǶWlQ��߁f�h��`� ҽ䶟R䯔0�	Uú�0U���2飼	KR��+BA!7���s�t?��Y:�eE2����/���/.�Q8����MG6�o���!A%F���.�ٝ\�p�k�gxˈ��8���:	q�Bh@_D�C�y�]s[��'>SK��K��Yϋ�aV�����R�D\��a����
�0��n�F\���l��yh�y���f���)a2,�un@ҌG69,��nn����k��Ԡ�ټ��o�B�`^?_�0L��pu��jE��-�qդ�r����kj<�����J�"�` �^l��>4�?�f��AʕZ��;��Tt�7e���M�R>W�`��i���;ǉ�4:t$���[�G_J��2S��`��<��9��Sb��Z�����~�D�d,������*�Å��~g�����QB2$8Cb�SJS���8H��	F�PavA���T����u�>ϗ)�V!UƔs?�\��/��oa����d��o
Rh]��6��kJBB�-����-��[�A=0!o�F�f$�vB����<�?�N��1Wt�P��y{\��ƥ*kwr���nt�JzO����1b��K͞��
(����튕Fϑ�C�NYI�7�nc��Ӄ5j�2 �>1PM!��f��DN"��|t��'F�����&cD��ʃ�pKIy76fW��=�:y��\�B��
Vv����68W+0�N,��Հ���i3���k�̉6�w#3�@��u>��j�-��������#U���9=>��a_����O>K�GД~׃*��s���h �߃~�>��p�oV��p'O��:d�ɞj@�w#L@�2���,�n4�+�R��O�U�������L���q([�R�ۍ�n��4��;}��kɅ2�)��x�}�^k�<���RUi��n����r.�y��PC��u_�IO+Y�l���"�q��+K`Mᥧ�
_����'�!���ex~fI+{����9jF��?MD*���1�����3�� ��a���C˗���k�B�f��t'(��S���'#ӧ��'P��%�e�W�c�}@�\5Э��sS:01�0I,�]i�q)�c���Gq-9!��x}�u�i��_����]�̱�
7�}�qOǜ� ��N|��4e�L�P@2XǝQ�w�Ƿiۘ_�B'В��0q)��5���0�=��8��@��F�~%"vH��ةѥ���h�I��菠�}j�S�Xћ�dݍp��88�e}�x���[�1��!���~+c`���Zg��4�~�x-�է�E;�Z�w7op!�^F��OP0�@D,	"�i���&�x��}I���AL+2�����@�n�~����/|���@q��]�N2@�K�������sB�gY}K�#�mI��R�\֏\� %��NHJ���&N��!���0C�ar92��?�Q��l��2�ˮQ��XE��n�ǩ��t�>�d3B�nSl�ނ��������zqWu�����KU/%ZV��I7�1�Z�(F@�k�T�oX���ȜA"���GX��O�yp}���H�t�!a�g��!]m)��F�۰�ݪ�6<��ߟϯ��n3��_��N'�����oG�g���-G�F�,��f�i�|�q@��}�Eo�1O��o,��QJ�m��?ms�������9���c�#k�g-��-#ŭ�L�����eX̼�D�9T�r@Z��.��/���L�:5Z��`��Ṙg��8G�7��R�K�[
�&�q��؂���L��Y�*E�L/>x1��r��G�"��
|��`-<��-}���:};� ����)
~Żߨ�)n.�����\�U ���}W�V-"U����ϑo��X�6�m�,����ѝP�+iT�:�m����Cl[�a��� ��}�m�j	`�M�t�*凼�t�\Ru-��R��Ö���t.���fG-��G�蹡{د�~�I9o�aE��yB	���I�L+=��G�[I�F�,�v�
S`�M]J�!;�7�@�w�c�rY7t�y� �$��T��}��Vc�E��ϗk}�%���`=Dc�_Qҟ��C���v��}���$¬�jI�~�(z ����"Po�<AN�*B��14Љ~�����qU�>6e����M�iO����/��M�Ә���u�^��]/g0e@d��8p��U�����Ϳ"�����̐�p
��X%��U�C��Se$Lj���p�O�*)������/�c{S_�AޝRZQ8	SZ���u�v7��@4�7$����%[ta����%��d�� L�f#f�^�W_#I0�J&+EQ`�໼�pN�5��-t�������
z�آ%h��b�M�,��ǩEQ�g��򗤚q�A�� 7�.��6ҹdN t�m�O3o�KT�-7�Q�~��V1m{2��I�a�xq_�KWǉ�1%ڀG�6r��c��N���j��*4��%�7A -��3�jE�:��^�����?��13!�����$Z�y�L������}��\�������������zaB�;����J3�ϳ*�g���(G�>Z
�?�
��(TX��Z�N!O�4�4[N��վ�����H���$l���:+j�T�8�){�Y$~莂�QF2ڧռ�� S0���7L��b�u�� �@ޫ2`ye}nHx��J���Q1�Vg^r%�G�䅘;�����@�SAF�:X�Fe1JQ�l �:�a��R�]~�t[�]W���A�J�!��ѐ�n�d�I��J�Qz�.=�	��Q �؏��Q���"�2/R�߹�90�%3�p�1����?��G�#r�����S"L`z���V+`�5l��v	>Sx+b]+�'*��?H���!�s+0��,A��F�&ϙĻeGn*D%Y