XlxV64EB    19ba     9c0�A�;��ʽ���v-ĹI����_���? /�ID��5"m��UN^�A��<��Y3�Ӆ����mwݏ�t��%%>�V�C��l�+9��%�Ub���@�.����e���ԊNn�Gߡh�b��Q�+�#"�t����O�R<+Isg�'�xz�j{E�g�^�Lg�R|Q'�HJ�#�n�]�i����]���=;�p-��|�B���
�1�j�L��]��-�c�G���+�����B;�fn������7�R�U�<��~��A��X��83+n9�Zr4E�+��w��">�OM�*!��Z@�ۋڥ�����~t���w�	l8k�&�YnO?�ܭ�A翋��?��@`Cn�!?�O@�I�_w����E1H���;SR�+�7���;��P�[�Aa���+3D,� #}�b<���W-ր�яܘ��@�R���)�V�L�u��M��]�}	Ҹ�>�D�L�QPh��'� �����'�0e�2v-9�Hlc��Qy���s�����~ni'�M�5�:��}x������������p�+NX�u,�-��rk�`	-�y&K��
�
N�R�t�4b�?��A�p�r��^�j~B]"������0�aα�d����z�+-�)����f�G�;���OդT�C��Z�\f�F+4	~x�h;;�1����������q��`"����)��l7��憣E�bdIJ���~GB�1;�L�'q̕$���a��b�9�[%�Xٹ*DP�\Ѯ������A�È�%�M}+"��pbO=!�*���a.����ƣ�@A�4�c{��ݐ�$�vw���Gс����]3�?s���v6mvT����PU� +�'���Ua������K^ȩ�0zH$�}x��hX��h�h�iXWf���)�P��f�I8�{@d\i3FbG��h��N��$\Br��"g�s@F�\���şa�k�M�b4Ø��GϿ� �'�1eGz�HN������3�8j6� �B^��A�=Fp܎�r�n�0%j�Ph�X@��sP#QC��H
N�y������M�]�-b��2��*����H��[��~��yA�����P��Cź���E-1,�:��W�&��}p(E�cc,`E�K=4ǧ�_&IT��n�u;��>��>c)�k��d�DHo�m(�|��>�B�A� �AG[g����q���Ha-�����P�r�K�Yx_)ωtD'&0�ߌ�L� ��f�x%�����jR�-_ w	q��,�
��P,�k�U����E��6n�����`P�����@k�/X���>���y�{0�iȘ��O��d)�O�����V��XЀ�\�`�w'�eD�h�Qb�f�z�m���K�}�Կ����i���W��Ƚ�Ӟ=cQ�C-6�W$96�Q�sy�rž��L�q,J�]���/O�,��)���җLh#o#�0Emмì*m���G� ,�ۄ���Cx�6�2z]�Փ��X�}�+"9z�����q{���r}ݪ��M ���ά[��>,�#�E�;3h�mkA�U$���Ǣ%��H#�86�:��>�抏h�갱��{�0�"F4�UI�(ϢX|M�{(D�P;% �}x�{�L]�_K�r#<b��^_q��W$/�O���i�8����w��gkb���V#�>P��#�;4�qٓ�b�_�X-/���=�kU�:�A�s���R2^Sm�P˒��)?��n�rO�����`3�1��~EO��eTFN�Ք��L�Jp�),G\�v���ۖ�U!�������u>��i�y⸄H�����I�/0����z@&��N$y��
�9��0�c<~�;��e^���l��D��B�qk�9A���s�q+�d�z@x����)Ȳ���b�/�����D���X�2���庉})�F������:�1�GH~�O�_�hS���d����Sk��n�|�,��\=�1�B����������O�V��6t�a=Z��$E����t���P74�h%E����ݔB[�!���X��`�J����x�ݿ<��ĳl��d	�/�T���9�
���g��Ѯ7��c@��'���ocY呕�7����-z\���q�H����݌�3δbl�W\�_j1ִ�Yxx	FIm=!(�F� T=Ξ��hd.+��:)�u9~��=,u\Q��)��l�|*8�괞Y��F}#���AN���#�s.kC��<���+:�Ǜ
�]k��A4ЗW�u ���e���}�hSG��{W�%J;�b��׺����(5�c�9�o�HI�x\�E�����G��>p�P쓿�bT�"��tH]}K�9��KaFXdo�ݷ�Lg���¾	�rOAbP�d�Ϳ��g##�\��È~�Zt���^tk�Ir�ԇӄ�����i��c8;�*�Vi��8��g}����}Dt:�i?ן��`_�R���1