XlxV64EB    5896    1450���pX�'(4N'ؐIU��?f��|��O�<=���w`������_H���>.+mT[�H�
6�biIVoA���#_ˠ~mu"vX��G$�Ȉ�O��������̴V[@�b!z��t:��	�]�൘l��[{��*�d$m.�jx]U��  S%K��Y���;]��WQ��[�צn�Q�'�R(��g7<E(FQA�2��)�=[:<
i�����%����� ^\t���ID�n/�����zYĊ���e-��C�TQ\��L���+:J�C�Hpф�Wd�[y2�<�p��T���2m6������b��3>�<%�JD3H��8��
T���/_�z2d=��V�9s�ić�;B����:��:��{^����"⑳�zu/2	$FL*���M�-!şy)ˊ|A�m.���F�[}�n/uت�?b��䶁dZ6��s�/�I�S�np���|Q�7^P�j���#h�U@��g_L��Yөu(	�t��y-F�2�pl ����ϰ���0e��ӈ�����Ti��Ś�$�$2t�}nI��=�.��|�Ѡ����i4�͸�%#��"N��Y�Ɋ��$C* ,��ѓa�ݴ椩�M�|
Ĺ�����I$�x����XI�E����V��V�d�>�*zz���-.7�v��P;�4>b��2M5R��Q,�������(�G�I����ҥ��n���"��(7,��H�c�Ikȑ*�Z��$���߰w�톭۴�y������Sژ���,϶��.��D�� �e;	̂N/�.�����$s�O��YF����S��J<'e�'��[��I��Sʐha�L�[X�����ߤ�oo�//
⧗c%������څAr���d#=f��ʉ���ؙz�Lpf���sgt�s!���pR�ӓM>6���h��X�K��a��+�e���0��x�{x-�]U�l;�	&��ʿ�~45H\K�j��F�w�NXEZI/��Az�Q$��J���C�VjCn#���##\�����	��G���e��2L/,\ͺk��J�����z��H3pdvx��,^��1�u|!�'����~�8*,���F�а�S3q�ն��&oءz?�����Dd�5��I�tYQ��=hҶJ�ڐ�y�r̅�j��y�����F���춫u��{ Fn[LRs�����'u����BX��%m`�ih1-���?-�ܼ	od�˞�QmlJjv���?a���kp�	�ٔ�U�t/�Y����`��u������ 䙺�=UKp�%�&C����)��C]�.j�2�r%rdΙڂ'ƍ]��Bu��!i,dL���4Vʋ�^ŧ
����V�ȃ.2Hc[��PQ�=���K"��a'Ս �Sˁ����n\k�U�����5��&UX4y��V��"�})T��(�ƣٔ}�~�i�mPD�j��ЃQ�4þ�m��&2ޜKFT��u���i���n�۾1��3N3u%���t��%WH��,�J����{_��sM�������f�a{�B�  >2Ҿŝ����c�`�t��,텏:��j�,�@���7��b5]�D'"��#z_*oIɚ!2�~Ikg�[8N?hQ>�{X>�;��O�GR̞�_�V�%r�T2t����,Iv����;��2��9|^��[�&�p��eđ'L5}��Ė��X�6ԟtU)�"r3 f��� �E�ʱ��ߞ)Ra�ʄ規�j[z���T�_ژT*�6�X=���F����P�p��O4���9\�؈�˅�D��_����~k��X�yh��b���tTc�1�&\�S:����\��ނ�18w�$�����sjӮ� ����<v�w�2E��qYȧ[J4A�e�Aq����>�r�w/��SX屓�1����t5��]�9c��jj�H4��9H�/Zj�������B��� >Q� ��#��Q�s�iP�P3��$��B�{�����������y������`PRp?`���p  40$Dm����;pV�M��fH�'�rU�*܇,ؐ���1�~����_� ��]~�z(�۰SF���x�{VrG>yGŨ|(��De�evQy��y����y����`N�Y]*=Lt��ʜP;�>�GU���0�u����V��m�	؟��:*�d�)�
�߄�3`/jv������G�P��Ss�{i�����RX�_}e].��}���|�S�/���~#��I	����5�>z2����?j���R��7�w��݂|{Z{ޥ	�qގ̤?��b͕q\��dяU�일�Ѹlp������*���P�6�ʖ����%��/��B���Q�U��\�B�����܅�`�l��0�VMds��שz���G��GV�R(0���M�X�c�������^���GǺT]4�f�C�������2bqlM���q]�"��A��ckN|֗,�w"T�n����e��P�HyV�N����^n�귡�p��T}�$1�:E�Ա��XV����|�6e�`�RP�o �1��1Xb$���W��n��^I����,܎�l.U)������lQj��:AC%g�?QH�j�T��>#�[�H���Ò��5�O�q����cW0Al�NH�&�%-�;���
��×]`f���T�:�*�/Z�w٩V��g�w�"\��'�k�7(� ɰ��Ԃ�#o��|��h���ܮ7"�(^c��jʃFB�f?�����~U�$�� ����-ѿ�"ٽ��'�m�;8�i�Ł�Ւ�4
Z�.~0-韍�BNX�p�p�<<�v;R;�S��L_��������b�x��K�X���0qV;5�s�̆�X�G�|AH� ����j�l��xlk�"Z��x~jǤ��̅�F�\��rC���������d����hk b$�q`��v���"8F�7��LԚ��)-h~$ދv��$�ZFw|:wS)+���Y�����f���v�Ch�-�+�����<�_���yؖ�"��E1GW��Vy��ǭ�8B��Tu�w�����Uܮs�lpKpП��"�6W�6Eb?!x�݇�JɸY>�YB��R�d�t�<A[}{{�i�y�菂%=s{�"ͣ�����.���+Ň��(���%��T�&�O�	�F<�jTq�br�y�Y��̔
�u!�&I�?�Q\��j����a��"�A	�.^���V���C�)��N���~ۚɶ�'��������:ń��w�Y��:����M�~}��$�s%�s�li�y�%ν��K-�
/��2x\y��Q�Z�x�z^Z��!�Uvi�飥�X���G�� ��g��DKMc��w_����X'���l_�y���A�AT���K"Y}��bh���QA�P�����1�25�7��D�e����d�Z\���Y�B-���ܮ��y���
�Z�V�n->��;u4˶�D�~���g!-�K����l��u�Y��u��E�޳{x��3NV�� �"���&|͞�͊R�h�ִ%u\R}�n��i����5�'��.������E�h���� v�g#q~������
����?��=2ɆwAD�Z��wM����/��/���e������rm�,�J��U-�����&G��@�"������;�o{����P[K^��^�w���7D�۝��P��`��.��b�V�OA�&��Q�~�����R��AGŌ���m�P@q�˾Y���MZtp:�8��*���hM��jo ���j�]s��V���d���`��OXdQ�vsE�ӨT���Zgb*�`�ӔK�������s�2H�#/�FL�EMM�K(�B!�2�b����@��4�)�E ɱ��~��9�b�*y��m����H{�a7;g`�q�O��2_�*<c$F+���B ohO���8o��^�O�>UЃ������ԃ�m�1�h^�����`����@�c��H6
ȗ��чq��Y��j�H&>�d�~���7j����O��{â3�ϐ]�x �(�,n�^Ҕ#���	=�5v�BpN����R�:���<Jtl%�\��V��^էF���D��0��C~���,�V�|9)��OR������7&)�?G�����hf�E�<��,i���V��=PC>��(�0W]&-�\^1x���󍥹M��7�CJ�����;�F3�ڼٲp$e��
8���� ܓ7�����Ss�C,J��fخ�jv\A�ٞ������tD���,���b	̶=�蔰����6�^cr��QD��Ǘ��[�!����a�\�z*\p��>o�I���𸆫��B��>�9XU*O�����;G'3��#3�Q��U,ۄ� m:�'5���j�2rw�_�\�CcN�Qg�xՊ�NN-�Bv�uG�\��"ֹa఍]CS���ܖ���mE��͏�j���>�3W��`*x<|��B������
��@d�m���5�H�MYSo� �6"�RZ�҇����`xo܀��ry]c3�����@��jH8N��TO!�Aw�0��A�l�);�v��,�,� �?&�O�i^#C�����U�$2�Z�g���7X-(��+����{��e���^fV6�8�E�������m��V���a@�.��AǾ������^=2��jy��N��O���-Z��vC�m0 }Eh� �G�~��������}PRJ��qX	N��*�rjQ�.���Z������?��5荭+�h�n� �Dѭ�v�p�ak,�ix��&�.,b����l�jT���z���(�1���qc$ ��]&�x6��m)��v @~�={BT<���r~��Ɍ)j�8Y��x�ڸ�v"���X8�1�U�������H�`�H �K�/U��׽�[X��[]�'�n�EX�u�U�'^��湐��?��n���)7W].�0�`�u��[�ҕ���	���u?K��O}{�p O9CY�wPև���ɿ{��LQ8���M<'>�1�gW��݇ly�r�p���B�=V��.-�@U7t�DC=�*��Gw��՞���nc ���!���o��p���K���HK3�B��^m� s!�C������0
Tv�M\2