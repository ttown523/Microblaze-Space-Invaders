XlxV64EB    2283     b10HcxF �]\5Bm)��(^]\?� (���RL[ ���(�>6_)SS$��J��Q	���*��!|���e۾�F�!���aM:.g�:}T�����$���Ɋ|�)��j9�j[�u'l��>-Up��v1z�ܾ��+�M�;��d��YE�śz=#�PR,�Z�Xb(��ߙ/x�ڼ�,ps D�5�*����@1������k����Ƒ2��͆~����F6���G*&������'�	P?5	AdF����-{�쒯�J�1�'>�j��ɦ%ɝ��u���:��๫k��
�l��'�� �aj
) �-�f�jja�K�� �� �ye���/�]�M��^2"�׿O	n���ê����IH����� �Vz�������g�8N,��(��ifAĨh�s.�'�1}�$��G}[]ҭ�5����l��s�� R���ᗒ<�ַ$��<�m��v�.��A�h��r���M��	�)��6���#'����,���Ł��-�n/M��_,�uD���.~�J}8Fܹ�`ڜ+��� �K��'���b��I�<-a��>\$4h]�t��<�*R�$����՞�c�#��|����)����!=��FZ�]�I��8~�C�y�����Z�5]	�w�ҘT�����xDk.�g�?ɂ.�̔�`X�k��mn���R�/m�K�v�~� �A;��W�g1�I>q�P�Z^�����Q\W�fO�Gy�Gw����=|�R�?]De��,��6i� /��v,LE^]�R[�;L��k�� s�������'[�K���
��[���(
3
�k+���t�=�� H1�7_bѯ^7��?�D�U��W��Uch�r�t((t�l�9[�n��V�o�Ti��f�͠�J�N���R%�[�}��r �3߂�.d��-�����.B�K���<����±���^����0�>2������\�AL���2G��I�7����D��ɟ�|�J��e�{�e�F=�	��|c�	��j[ �7��X\�d[H��cԞ�̖���:�����w�#�cf�����(����P��8��.�N�ߔ{����"�����8���a0P0�g�b��3`Ȇ���ӷ�G�,�j%6i~����П�:)����ȶ�#�&$|�O8Y63B8xNg�U+�Ow��l�D���7&����b�n|���c��\��h��Ί���߳�ʰ��}$Ӷ���z���!4�ٗ�	��n�#˰��Cc��[2���U�������8@�`Wz���*"^����ś��٩Ӷ����lIxH5N��Ā�c�w��0�v�x&Ә�}���¿rD=�k��BM����a~�0�m�)|w�̢�t�7^=�Lg�L�X`�[���u<��P�������S
��!�X���h6��X&؁w���%��ɚ1�5 ���o�!8�Z��f������,jrq8�ͅ/esFҨBD��j�>��*%�/[��XmR<*ٺ���5Mr�~΢E,�Q�J%���b�����%hn�+֒�$O�+�ͳ`8; Ə�^� ��o2���͓���,���8n�Y�K�F{1�ޅH�*��'����T����Y=������0�� �PVc�T�'��67^1�bP˿sΖ����r��65�zsʊ�v���k,��lE" ��2F[S�Nd�Z�\Y��wbFp� ����X8�&�|D����zN�k�W�A���5�r>ȑH࢛@RH��ߪ�D"�R�XZfݶ_�U~!��l�H��X���9�~�B!?�����w1�>�/w�7�92t׭k��y�Ϗ�0���݈`��9���g@�<���]��F����C�7õ}v&Dt}�$Ko�u(4�;�k�[�+u}���(�C�ڿC{v����`����mKp��BD��Jox2���l��f(��@W��Wj��~-S*Z�i�oI�,�����)<�a�0����SÁje��1��������w�ja��彻s��x��/�h� ��F �%C3���[dF 7��9.k߿G~W�%��|��
p�r�0R�e�?$
�l�7�k�g�A�<�?�)[���������������+9���E����x�슺�*�l6������"��}����^�o�<��`e�p���[����	�4j��٫�砠m�r?��k���k�$o�XA,����lM�Y�:SnU��%��Z9�d�}�Z��-����01!�OZ�����m	��QOz�v`��(�XM<O ��(��#C@���;�-�y����vC�߇��r�"i����4W2֗��&2@��(��M���w��7*��0���F����5�-J�J�Q��Q�YZ��nv..֟�O�����hP�;��9�X��-=t������Ǔ��\�+�-pY}�������Ke�� A}����C�,��L�u�#'�D�}��Ǌ��0��l£���bh���Y
f ��6<�=k�n�Tp��T f��bIE9�i[�S��^՛��E��(��ߑŉZ���D'F"�oZ�	�[�<2�o�����Z�\ˁ?v�n�i��ϫ;A�w���QmRс�cEb{��WC�����X��;�B��_�*;KN��&�ٮ��	���x��F�"B:ޯ	��H@�Y�L4�4����A����i�2z֌��fv�
�up�)�H�]�E`��/�0�l�oߎ�~b��0�.��(�l�y���J-O�9*��L'$����>.xo�%�t	�1�Ma�u|q��bŐ�*�Ǯ�^X�