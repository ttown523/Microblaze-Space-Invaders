XlxV64EB    fa00    2390+М��/0ȵP���p=k]6Q�]�D�?(��0t�o���=�-��>j|珸IU-.��i��e�gbN(�:��
�y&��|4�_=0#}�,�fnXo��CWI��E��a����^v!]�Z;;ޮ�5dB�kNe�:#��?��_�H"%U�MV8��K/ʘǍH��tӀ-�+5�e��~�"��f�#P��0�0�SnE�S�FYT߲|b���N-V��=�a�N���T/G�Nwŵ_)  �g��� ;��hS%��P�v��b�i"hvݚc��ۘ@ڌ��з�����a��Gj��S�o���1
�ӳݖ�q`�ʆ��Zbm/�&ω���8�|�8�*�lRQa��CX���土��&�ٙHF�y��"�IN��j�P����bX���\M�M���[�9�1a ^��6�x��&����i��h�i0+LT"�i#q)Ņ��zmjB2e+�S��mi�_N'�+�!$L�%x/�\w��_< c�,FO`f����܍��o�Ǵ��7J2/�B<�=���<�5 ��5��܇1V�JrwT���A9�F@���c�T�mdk�A�t���(�4w�n�W�����Y}M2�"|���#�-pڮW���j�۽t�LA��4����͎PH��Ix&�pQ�y�'���G�`\@?	�=!�B�F���M��� 9߷�Ԛ�
�5���G��.`fUI�pz�i�<?�3����}�R���*��А��+-�߁⃡@ ��Ϭs��"g�v>�Cӕ�،�]�H/���nMD����\2�������F��Ҥ��O<�lB��)���m�n���'�i ���6/cn3s}�ѕ*g��=�����"%{�J҈��rB�FU�q�����~W̔$���b���K�m�d]��^"���J7?��6V�R��>��g{`�Y�l.Gt��n�6J���&��4��V>�����TJ̑NL��˩�{4z������Z�$�A�"�:Yp!>'���?�"*[E�q�M��S'�3��l��Rp���\��=�d�]*�����i��5�ev؆&G_�Ξ���Sşw�����;�a8�~EF-�0T�.ވ;��3�k��{`&�K0y��$�<
^���
U�c"��)��:T~j?.�1��$yk�@*X�9�z�u�|1	Y��d�]u�eA��ʫڣ ��3��n��&��1����U*�%�����b��ҍ.Q�_����\����W�k[�;�5� ���)�k����Z��ύ��\/^�F�dv�N�Fd�T((-�6��&�/��C�d�heo��
-�TBO�e����#��8݅}�Jh�q�5��L�ȡ���Xc���,F;9!�(M�@$j�(͖O.�r��!�	�$pf�}��%��ZGR�_bx������=��o7g$3}-����N�#d�>����GCC����݁ߎq$)����ņ��w�}�s�|��r���m�=�����7����Ԋ^�Զ�F�7���$+ru��RE�����X����r�ɒ�l��k$��k��^w�7X�(��P���l�,�o�,�٢���q�u`F��EH�Yާf;��,���Kl��,�ߙ֭y.D�]�O��Ut�>�o�au�c:���t�AO1�;p�v~L���q�����P�������si�*yRY��&v��Q_?	e9T�DR7��mE(B�c��y�3>�\��{k>��쥕xu6�S��QBƙ' 'И4����<�7��͝٫e%�K�
�},��,���c����K��ya7��.�9���ύND�'�WDQ,@~�"��Ta}��1��6�>����u:�.N.,Ԫ'�0؊�BJ�����#�o�u2��(ݩ^�Y��tQ�E�hlh����F���ьOyĹ2�|���G O�!;������9 �ay��s»rx9�Sn�iȂ��f���<�,�l9
a�k��|?�����}��n�œ��x(c� �l�:��%|�Y�LH��,J�3a'=��X������d �	!��G50��~�_��/�!B�08|qD�+�XAe`�_�P �Q|)"��C���)�b
uys�H�Z�12��m}M��н���Ņ��pʠ���w'���g-*�,f���;jG����K���m�0�|��]��Z�%�!��;��t�UT�<,YS��r��Y��p+�.�IX�?4[�َV�����/L���5is)T"��.c!)NW4w9j�ߩl-\_����i�GE�5����ŻL#���f����	�ZT��<���"�"������	.
��]�	�9��5R"i9���jJ��y$[�q���4kgö|{y����]����~��;������.�&�E,�t�@މ�ai�Ť�qT�$��]��s�K�n�ʍ���j��M��Dc� \H�J�d�'k&�;��\x�:6���2���"��+ɮ"��8�+V� �k��Z������`f|�%�Lr7;�Y�h�l��k]��a�����n�D���>�w�zZ�]���^[�j����\��A�r$:�Y.��탞�۳v}�p�pw��W�:'貨qB�e�&�6�%D����j���SQ�p%�_�m�L0�EO��L��1g�(Fi�Lk�J��y�Dq����3��L���{GEM�6ph��1��Sf���*&L���9���g���.����.�=����!Q@����*��i��Q�G���.�	]y~��JX�(T���� M�ww ���l��Ac�<��)*	�DP*���1I{V�j�����-���R1�F1*)y�+��W? u��^s\�a��x9Z��
0���)K�
	��;f�rck�y{I�G�`��2UUn�:l���6�h�0Qy:Ƿ����*�q�hb1bߵ�w�BC
6�C��|�Zf8�2Ќ�Z�����;8�%Ç8W�k��?�+8 �̚�zrp{�DK�+��VI���c�&'�8]E�Y�u�iЎ==�H_Ջ�pD�82�a�~����_P�E��i�{f���kª[�MC�ϐ�
�@�<ho��D>����ށ��[a�]
?Eg>2��z}�drA
�R�ٛ�DԒ��Y����p@p�M���Hj��ʎ��b�jg�ȋ�MS�U�&R(��`�Qp��Z��u}�<����Ҽ��H�oDR$
xx�0�Vh������d�Р��`v�)�2mS:dM;]C��v�8>rQR�T�<5���W1M^>��u0i�����.�͇	?�$�8?��(f�-}��!�ZXN-��jb��EeH�6��xz!t�S�5�e휇	(9�����q�PX��K����_U3����`N�u�Qt;&����L�@�P}�O�by��,�S�;�|�M��	�s-��+��h#>X���N_>a���#�n�/�3��Z��E-����癸qΦ6�KDrL�5L����m��9�W���/u>�@�̳k�l\;�״���]v6)�[�$��al^��S'8��n,��ȇ6�:���PF���ˏ��}�a��?I�a��
�����K������_\r�0���8�S���v>�h����5���{O�����X�Gp�2�1(�hP�A����z��k�eW!~Kp=o6�柮{nn<ntF��?��d5í.f���Ω�ZΔ�-��&}�#�j�SX[SX�>�阝#���N��o5��W+�г��ux�.o���P��9å��ID4�1G�D��F1)]X�`�B]s�%@���r.�ՒX�x�l�}�Q�qN	�}
��?{ͣ��L�����!�<,$�U�#9�� �s�l�4�SR#Ş����fn@���X��ݹM��
���.$��T�zv�L|�U.�'+F> �S��C���~�RD���!��us��y\��eE3���*�-�2��AOk�l=�5�p�9�D�뫱���Ç��rY�(�˟�5'�����h��cm���v�hV��Ȫv|���&Jq���C}��A��Z�g�q�;xa �F�G=�
�;����f��`�������%���ß?��ט��mݹ��'/���:'������oJKOnt��Z��=4k84�.�G�H�:�mm��c��4�"�;ɮ�n��rղ��l N���ќȐ�s��,�ߵ>�����egPBAќ��E����tr=ޓ3-x}�����<Y|�;芛0�E�����	�W QJ�i��M]����}�ˇz{d��{]���E2�����bF�顓]�P���=��,�ͣ�0?�3e*2��[w�#��� lnu���~��,7�� ���;Oݼ�m���t�K��h�Ɨ��3�� i܏S6�\�����tԿ�����L.=��XE�#jO��#nHE�>F���0.�j�P�"kxDuԝs�o��,�g�ܼ.�ƙ��v��ֻ�S�I�/�*(���h��̝%����N ���-Ēq���w�ᇋ�N?1�2�`R���h�G
���q�J1��Rɫ���������%$s;���C};��t�rP�0z3_��X~N��bc�8E� �4�Z0�KA���2��d�������`���B�:�R1W� K����<͊"��@>���ꚓ�d`)Q�=m�Q�F��=�ӏ*�	�*�+�7a�0�.ڣ_�bU�ȫ��g�pfK���@H��y�F�(3��¤;7�:�n�����#��j�M��=K-t����'�ߗڤ�F��`+Q��`~���b�~����J��d�d��;=�ݞ�	����']�b��TO��zd�Q�J�uN�#>�W�!}��j\�ڗ:q\��oC� 6� i�+gPX4�&N�Q�/��R�CD˻?������e��{X��r9���a7��prO+!��q�&{ΨOn!��
�d�A�7pL�6r�.S�8�&s��	(�y�Q6��[$W>����n��������`�V����W8+FG��K�		לIY�����[Xh)�!��W���"VT)��U�t�]-�7k�����B�^�PKxe&�M�]+@iu���|��@D�^G��!Bn@*<}~x�� ��S�B�+9�R���i�alm|�!g��� 8��(����_�*_b��R<-�dAC:zg�籋Tڗ�{�&�a,�l�����>ei�ܩ��dG���S �i��~K��>N���	�[_k�upmj�Z�4�&"{4��^|�R��2�����X�I��6�����y�;��Z���È���ȷ� �V3]���:FGǘ��A��nqub�^�� �m�hV�.�6t�������1���]���ZÏ�������+�
�c�7�[rc�3[�&�Q�<pu��	�ٴ�j%��7���_D)�Mn8��K�sc�2>3@Ҡ�hĬ�5`�d�R��D*阨�,���L~=�X�����'�|�Q�0�"�3�etv��E,qK8 G�4� ���I��&��(y(%�j+_
�����&����X\��W7FhM@��A^�AEf�i2�������.�;�"�ċT�U��xz��jW�Es��>2���g�nh@I+F��hV�]�9*"s��b����P$y$
SA��>/���x}��Uyb��M�P�5��Z} �x3��,����5�A!�P|��J�%S�a�s�҄���S����/�~2�Ȏm�5%@��x���t��]�����fXqZ����lrֿQ�d����b�K���1�P�P_M�]�Яa}�B!��SGLUUf�"(�0�	�ͧݜ�$��-�8r7֍��xG��DʋSM���w-�W)5PcY!;,�kF��kp��m�?EEa_}�%o	f��C �\��}M �_�����ǅg�}�4滚�M��F��Tv)N����hq_)�,ͳ�����v��Է���R^$-�@�@�И��t�UN� ���GG���yW7�/��3���k-�)�M*����A�M��9�֔c^�.�Tx��+���h(v����Cc#�gx6T��Z�*�9d5Iu�2yQ%aDT���(�W��1�W���0d�j��q���k˜�?�o�0�>��k�F%�� �#!E2�Y�e?+� ߹U�t�� �iq̨�R�?L]5�a�v:���}���;c�X=⤱�m�]Br��P:M�S���ίgW<O$Y�
l��t�ʦ���R4y��̳p7�R���@��O�[�,>�r&P�C��bKmOoe;ЫĐ�zʭ�䎀�J�M��'�i�
"��Y"����2��G.�&i��juv8�t�L�Gd������{ A'S��d�����HT\8�G�c����ҽa�/-J���+)!0~���s�Gv?V7���-l�Ӌ'���DjO�M����>4��ڂ�2��M@������y����5�a�縸�7 WX�t�9_-��V���D��^a�Pr�@�tRD��/�q�{����4���L��ڠ�����C����"n�T�+)�"� ����]h�����c�ѳb<��JL@>�{����2�A�"�0-n��!�q�{�ʣ|xфa1Qtj�����e
�+g�
t��LI�$�x��S@������
�D��˰� 5�<�]Vy��㎜�|���}�� � yG�F���T��ȅ����k�3�̩BoFIc=:�I�nF��.��u��*�Xv$�O� �f����>-ZǸ-������������t��O��Ӄ�b��#�P��<��y2Lk�P>f�E�V򿥙�Ax�����3�9[J����)P�W9_�(�ؐ����X:�^���9��H�Y !]?���>�D.���ނ˳��^�ϳ�Z���w�-��ؙ<�`�3���F�����UZ/��dFfݓG��h��(���Kf^Ee�֗��'$���A�Y��E�_׆���!�F�`<�[��"�|fj',���Xn��\n=2��{���Z���U�\������cRPcABX�{�"Ii�Pu�*q+��_���
B�&.Tp���P�]{SA��7?�iBY�����^�rf��<��4����|�P��@Nk���*���@��l ��)If�!��GƯk��;�1�����
��pY�p��H�7��L���V$����<*+�$�"z���5�9�J��S	�ŷ���մ(3��ē���^BSg��/p5�� ��.W���ܳ*f_��N���-��.�f�-.;W�o��[���z9H?V�ex0h�yL����=K����k�����Y����Ӆ���� IY�=U^���a�w�б���zpWJ�ܔ�`�/���|ǂ[M�t�?X` ��Ȩ�6��#�L%>LK����!��2����vȔl�5#NA$�e[�2�8��:���,߿�,$ڷ8؁�@7��fS� N̴aQ%��A�L%(���1�d�
$�6w8��lC�iS%�����)�ڂƏ=�d��;�t{���}0�YP�`��n�;��3s$���Y��.P,�9#h�e�?79Ep�0���/�#��S���e͗8.4B`q�w�Pq�BVX���0��n��r+�{��x�|@K�~�A琤��k�d{�ɝ+S�t{�'���J(�OO���p��?`�;|B��bJ�0��J_�08���������I\�������Z%�`QWb0ڍ���H�P�V��+`�p�<U�c��<]�aC�H��{��A���2Ok���\fm<3`R��L�2�������װ��zڰo �u��p`�p9�𐣄������a��J�R^���?�'����3�U�k8u��SII��4�O�jy����vP�qC��}�4)�~E�U�j�p����;�P�	Mrb�GIY�P�	7��!����W�pC܍rwj�ZH5)L&��'����*A��i��lի`<[_:k&y9�H����u�Ő'y�ד�#	|��7<:�ѲD��3q��}��U9)e(Zp�j�Fcn�sv��c�f����;u�b�\M*2@`�眵�-Ϯ�7"ft�B���a��_�rDj`���Πv���OQ?[R�˓B@�si
����ֆ�Yj���$���)|�{*7���}�=��&�O@�g��DӢˡE�m�ܵ�������+��Y��gGg�oi$u�]��OqP�����:$��.�U�|�f�pm��,d̀`�8���zF!��1�@�=k������܈,A��J5�#���N��XQ�1�3U�-�:>�X��~��so=��ۈM�7��l������ߗ�`����0�9��[�
Ĥ��H� ��x�Y��E�w�܏�INI�ȍS˜-|�	O�<) �oA�k�Ψ �/�Ɠ�������%�qn1=ti�嵓7r���" �|��J��р�Q�����$�%�R��p�%�P��Iiw�Ԋ�	*
��$�ox��!�%�"���܀zQM(7��O��mO��joJiº���>4\)?2��%簹�v<�m^A���-�PiYU�K��ٷ45���X~X���r�_p�>�)<8,�=�����Kjh����,���뢷׀g�5bL�Rm��}R��>*�[5W�v��sԸ���3�j��L}Z�9m����[�d.�\	C�i����VH��)���������RDJ�M�߁�,���-Cp��n�#b:M�H�� h7��q2��>Zs
H&���)�kQ/n2�����D�. �I�X2�{���G���.J>U���m�/��X\.�Ĝ���������&��2���Ԋב����k!kJ�(.�ۗ��TX:���R��S���|y(��N6�'������2�	�5G��w��Cn���C�9i�f�h�WϏ��u6V�(����|�;q����oM]"�l�a�1��B��4L-�ֿ�JĆ��\�/
��y�t�g穑^��i��������m�M�h�0��d ?�ג�+� 2�[hӌN�żv� ?�c�N�b�pR�k�2XlxV64EB    fa00    2600{���-��ʔ��9���O��/?�94����Y��$foC`�'Δ_��:�#�!:"o�,'�`� ���T>)gc�Hi �UWT&�n&v�*�7z�g"BO�d�,���\m!�È��J�o��M\�j[����?�8�)�2�F��Z�=�[�3�`)�2.�#�VZާ��o�O�о�\>H�K�٫����b_�	X��Y��:6&�=�u� 7d&s�!��w�u�����}j������^u�\�a*�\�Fe���!�>�8t�%폹��̹"�T����p&,�e��������u�L��F�X���7�u�9�#�R)ņ����>]�f.�I���R�CgU��B/&L��7܎Y��.�6�w7tN��SsJΊ����ǻ���3�Vü����.:>o���}��/0�C��Gp�ҜeC7;�����H8��f^���������l�D��~�J�_0x���X�"�6Q�sY[��#~1������
�#�����I��p �I�v�v�3+��"�>�5�Ӌ��,�Fr*��U�GZ^�O�te+���x�I�A�/�5 �dz�A��:t:q^Ü�.Z2M��hW�{�����!��K#V�$RD?���>��e�:@��qM
����TT���:�Z���\T��.�<0���������D��^��8w~�$�i�g1�i�]�{���FI�3� ���V�U���L&�F��
�u�kZq���ySO82֒C7]Q3@�#QQ�LFf����<��o<9�co8�1��{�:Y^(�q[iK��(f�yN=���qqb~�$G�-�Af��0`fU���	�dYͦ'2B��Q��hUo�Ӿߋ_={@�e�dQ�+�17��<���z��rEz,�A��9��"��4�}���l��uk��S߱���H XFeԖ��"���N�����{�\��)�s3ھq��j���A�<.�����Ջ�E���S/[a�}e�X���m���S�=�A��4c����uκ�7jP���G�8'P��ʴ�3�]�m��g��A��Q�>���kRr讁�/"��/Ŷ�Pro�iW���`��[����l�K�����.;4h#Ȟ�
PFyC甃o����o3�c��S�Lӛ�-����B�� ,̳�U����9��iԜ�� �&�	�x��'qaҤ^�I�j�:s�	���RA*	�^��Sj��Ѯ�7Fi p	��H7����
��/Ԃ`{ӛ�5 ����P��稡/q�{ܚ���k&���z��H!"��&$r�=}�;^H� ��0�ƼK�*���
�� oJ����ª�@�ڙީ@'����>�M9�B	�����L���FK�r�}����meI�.�0���@��A]nt�:����w�g��A9����(:AEW����-�����B(�<����f����*9ťN�-ʰ����e��ْvXD�a�@ nm�(	�N��F<
����-�0BK8<r�V�������P̩�Tf8 8{�����Y
Ď^��l�˫��K�NԦ$�?�'�|��j4����=%���v�/��6�f����r-
4�j~���8���ѫ��ڏ��yo�t�������x� %7��);�]N+�[�sľ-SG�>Z�U:S\r�{9��>���(�3rH\ɚ���h/�����`u��h�9v#�gI�_����J�,f��*��YQ�����P����e�S-v��}C՜�`J��D�΄��7�e��y!0�ɑ����
v-�m�� �lbS�*�g7�_6������,��_J��&���sV�&kr������� ��ʫL����"(����L~G�^��*Ql�}�H{�����,S#�Å�t,�|���\E~��N���~W{�3�/���/ӟ�:�d�'`a1�Nʩ�)>J��4*�1W=���5�hX�d��펕��!�:�mH�Kh��
+4���������-����G�#'���~���;�r��,�\矯E�,i�����S%���r֣vo��Tn�J���n�N�����L����!����k���T�
��{�;9^���߿��cN�w�j�)���\���ߵl8��O��N�9o�Ja�D������Q��/���fH`�4 B��o�;j���� %���7t����9�]������X��r��V�*�f�����٭~f��&�Zf���Ԫ�L���6��#�b���ƾ�vnpY�<�Y�|����ݥ�4(��c��}r�W�M6� �����G�Z����8�Wc;9	�b�A��C�wb��7�m��X�*I��$"S$�������T�x�V�q����Wc���p��z��Ş�l�XXӳ� �����<�'L�d�Ԡ'ΤT��%ZV�U�y"�>�C2�d�6dw|X�-�G*dqx�.E"�_(�g�M����8�'��4��j�̘S5�#�t3#P
<�I�r��J���%����`4e�_�y/�����G�V�,��ҝ1��f�I��N��r	�d���������+*��CI�k6�b�i��P��J��ж.�d|�G���Wrn����L����^��{j��^��X��+(�,��Lw�S�ŭ���=�\�Q����jH�7���t,��(.K���A`������"�l� 6` �LZ��o��}1Ms�x`���raގ��!&m��/E�r�~`A �V{�\��,��2�9=v�Ȑ[���M7�y�X��p��%"	U'qŵ��iP��j�ُ `�{[[�9F�������KV�Η&������o@�Ov8W)S�Km�Q�^��B�N���"~�V�SNH�P!�oʵ����2�R�X¤�a�*�JBe|��	�,�- +��@���S2f˨�����ޮ�.��i�SDi�Z~��x�n�%B>��*�b�}�,���R4E
��+�0	B��Ԟ%+֭�%v�CTl�@�b�#�]�w�+I>���M^�CwtJ��n��� 9�����a�F3�����7���\ �S�*��u����[�i٭�'A����?y���1��d/=f湖z�z�5��� }[�P@���5J�c����zʀ+|�p�Է�VS[?m{���4��\ O�}���Q�JgH��R̋:�w�C0�G�lf�t�v_o�6,�{���#���5k�
��RE[�˕���()�e�@��5F,/�bР�n00��݄���}~x�-��Ɩ�i�90��z��=p�}��\.���e���4�q�]����y��B��޺xwbfa��Hgc��ؓh3(�!9W�I2n.N��g���$˭/]�Q�nr2o����A���`��(*9����_�LO�8a����U�״�x"�M��K�[B��-��q�_{|{��t�rJK�8!�s�3��"P��,�=�D~ePQ��^<˵��K=PPw���{�/:Ϗ��ó�W���Ȃ�=Q��W��\��-A�ͼ���Ip!�7�7�DNb��Dv�Klpj���j�1�R{�MNc�K��i��bNr����nZ-H�Sxv�w��Z�}�[-RU�F!��f{�$v�+ϥ�I�B�NǬ���s3{�P�/��E�˘�_O�b��@�'��k6q�x@gE�s�*��q�k|��O��i\�p�}p�$5_��-��@|f~���-�F�2��EK
���� ��(�T�XUՅ�3܊;z#��a���,$�[�{i+$���n�D�2!-�Q��3��hc�(l��i��Y�&kR�خ^1������P,`ԇZ ?�:�7{�e��R�p/;d���#���j �\�)��
��ʢ�J�Z�7b�����5�B�6L��nƯt���q���	�k>A�{� ��NA�����{k"��1����(�����P���a�� �C�G�O��]9�s�&�Go�<���٬A� KЎ�rᏪ�c�d!�0x��Ot��L *�zZW'v��3����e�hvg0޼s\9�Ⱥ')Bap�[��Q�������٫�2әJ:&r�
���߭~bL������
fm.=}��+��7ϲЊn�]�-�;�VF]q8��~㣬���jB �|{dB{�"A���6Xi�$�.e+�p���GB �z�Z�Hۃacr��˰�����0�]���|���ҭ�vkS��n&��("�7d�{�P����=

��$W�L�P��T)4?�3Is��" G��e��-ewaU@������A�����Kw;���:{��>_��Ho�3L$[��-}�O��r@�9�	��}�]ş�e��p�����:$��^�*A�K_X� Ը�
;R����"l�Y菜�j���}j��d_�������G-�a��lhD��YuL�ƂB����^�e�ǀ�?�p��;�/+�CʷG�L6
�K�_�(Y�	��ۈ�H~�y��gh��2?[�����	�e�����y����h.D1���t]�HT����0��.n��A��T�����Ke�r�rR���,�
W䡸#�lt>�-�
u�ׅ��D�о}�#�$w��2O���u6��+ܮ���D�ϙv�[�6�q�Y���pF�������˖C�n�,8���Gȋ|�4 �>R�2E&0�;|Ui`uN�8���u��ͻ�_���_?,MBb~�~V'i�<�I�C�z�+p����r�<"��R!m��$pӽM��L�v6��W\"ʇm�H�J�`ޝ����2��Z=*[����Rs�]����̴���u�u��o��i���w�@�M�y�p_?{������a�N\_�;Ə��N?�������ߐ�4po"�0I�/!WM���f�|i��jT��4�& v�$b���q o��1�&5>�4�$���)>�����D�/P�R����Ɇ�\�>)\a�h��.l�Ky��$�⦁)�c��K��_~�5�{�y��}X�U��!�Wf6w�tiV�s}���L:L�HN����f�G�R;��x��s;ݎ��^b1w�۔g�ёXQ
�6a�,���Y� U�㞽���l�[�Om��{��+5N��G�d@���{�-���#�2�2�	�r<6ڈ� ��B��W�oEAv߷~��}hl���,�	�̐G����c�/k�;�w��M~��Y;8�u�1(�?��.��~�/~��@�ʗKY���X�u��U0t,���i=�������j*ϰ7e�Df����V�hX���F�3~d� Q/z��%  �TR}����7�ݧ��������8e¤ ��JR�@�JB�J��'�)|��ˇ��i5S\ep�'b 	57���7��ƹ�˃qcǔ�[���ѰVJ`.r�3q]dOy(x��;F�ߖ� �qBi�ĕ�n-��I���H,L2(��+�
.l� �RJ��t�6�q�0�V��H�\�g�+S����9<l2�S���6����b{Tz
�ͭ���]	��:}��\��y-61�x"���S�$��X���1s�bEKA�t���o�䁊��*��o���g�����e5�o쉹�a\�/OP����=�բ�rG�&�.��AIP��F��WoK�O�f��L��u�W��V�]צ�@�/�ߢ�K �H`S}�e4�́�ן��]�K
����d-�1Y� N	�ԙ��ҽ���ֿ�Q��5��f�V�r6Z��_��J����ÒgJh�,`�s

̫\�}Ηf<̂���ZR�q�ᚃ����#���Y/� ��_�\!�v_`�2��bݙ@�aMɸ����Ū�&�З�O���jY�+Z4��y#l%�Ä�ͩd���Q�nYW
����3���F�yV���m�F�ǻ�w�
����w�*_�Jm��
]���_�ǡ�lc�r�`�'�E(��^��EV���PD�{+bR�!��E�e)��jy>"��-�MX7l�'ծ�?9�=w��%oN�	�0��o��"��/��[�ǘhА2���.�4D�Ȫ�;}ë(�k��|Ѽɋ����2Pv��'`�aR
��ܝ:���c�O伙2���O){w���:K�!+��A�۹�ƒ�L� �@H��p��5�/�s��f�r5`i5\_?�A�	�N�e�W��O�`��v1?Xl凉�W��+�O�ԑJ�@���?U�:VҒ�w0�o� [:�u�?��u�ڌ�:��Zc@�V�v���XN�ء�Q��W%#'�4Ǳ)�r��P1�=���Iuϡ�%�Go~\�翚��M1�Oʢ�K��H�X��xzm)9Y%#	fx=�D�{�<�?I���	�с�<��6����B4�rh���;���d\}o�m�?ks�1�;��1��{�^^�I��� U�s��燉=Mo�r�J��]=b�'[��8�^�DgL�Z:<���"U�1>��&�e�=.�2�Ue���
�w��m��S����!쾴_��� �ӣ�r�D[��W���E*+7�h�>��Op/�xkDEX��'�LpIc663p�m��}C�K3̧!;�T���[����^��L�1������v��X� c'�Īі�ݯ�&DhDI�r.>���[�Ka�q�D���@���)���W�%���Ꚑ����aA�:�)�����IR�_�j3�}�2�Le"S���_r▿���:�94�/A�h�цzi�#=�I�7�{���vh��k���.Ue���V����l�̵o����Tl4h\����}3ܙ�,��TVd����"+Q�x�)�d��<h �0-!��Z=O53&��!���P[[^�&��00�hԇ����n(3jW�{�{�?,��`MV�g��j"������PL������T{@�$���F��WF�ދ�Y����E�Qgu�������{?I�̣~�1=���7���{�Z�&��3��������-!��v|������J����/+w�������ށ��ik��p�`����ߖ��(�n#XD^���`��#�d�@2���܇ z���6���O]�tgoFs�u��ex;:�16CDC�F沿K����z�Mn�ks�;��hV� g@Z��P�f,�t������+lX#���Ŵo�,��_���5�i{��mꀥz��=�k������4����iڔ���X��PV�4��e佗3T��q����qI9�|�����{�T�w� a5f�J��]�b��ۈ�:(��ˁ�C�z�PQ�vs�Wn������x����j���s�6�����.w?1����	6���u�Y�%�h�ozj���%�x�����ߚNC�z���i9�ٙ�U,ϛ<iv���4<��6jV����b,�%u�A4`ډ�0t=�Ma~b�d��+�$�wo�6��0U?GP�x0���f��h��i�,�B�f��Q���0�a�L�we�aD���x{?�	 �C>����� �TW��0�S�r��׻TJ	�aE�Q�c���^t�5N^S���謤%M�{v[*ߌ������ٽ>ܹ�mo�SMx��hU	������8M\���~�n-��nO��y���>��]�s�����o�$���z�i�[��;�ω�~�WӍemO�@a��bpx���^��LW����H!��8������~�=1���\�D�5���M��UO�o�o\
Q�ͥ�x�R�S�;q�L�����Az؂���
ڂВ�xg��h��<*ʙ�����G��]�ֽ��-i�����M�]��8Qa_C&�U�r#|p^�s�Ǚj��=���c��د��ҢkO�1˱�go�H�ϔ����F�����\,5�iYмjA�@<���`H7��]k��e��N4���<����ce������R&��h�
e2�i��N`S�l�tX�u
�BU�&R�9�SHT5C;ʙW6�ֶ[/r�q��j��Q������ ~��:5%=��؝P������{7C��yKC�͆��ڐ���("�B�T����O)b34�S���j*�`��wĘ&��j�p�]�L�̪�p��<�W��Û�G�e�}�� }ZMF�(����v�T<n���|�5�x/��1�	Mn�4��M?D�Җ&�@;�s�����},�x���쑬���#l��9�Ǯu���{�$���W��@LP�.]���3� m�%]Y�� �VRO��M~��=o�+�b#��b��1���ZMz/��<Ӛ�T��z��r]�7y�k9>Ԏ�����hQ�Ք������ʑ�M%q��\X.��0JQ��w�������t+���M����@Խ��C�HQ�.��)���|5���ֵY�Ww�u�xf��-�#/\cc��1X�f=�󵐷<PK���;�;;es�)	����ٰ�P:ß�eTw��O0:�gٗO8-�&�
DT�4��I�ײ�����HϷ���R��4����?�� <y�/�?x�0�Ȥ�M���H�������bH(G�6 �h9�������V���h�as$�U������A9_x�@k�Y���l�S�$��t��O�0��'�֬�(���_y���E��(.��E�K�- �~�����.P�uj��:��z��,���O��(�}�<܂�(Mv��d��N�!����m��F�d�5�\<��$� �:^� eO�a7:��^��%z~úYJ��j�s�Q���)�摐P��sBP�9�6j�<�dAsˮF~��J�[��5�ʥY>︇�D�i�=���k ��ӭ�J,�B����b�l'�¥��􊃸<H�"��Ёb��i�}������*
���umq���^I-\
�zz筮��S�ϲiňj |�cu��+Q�t�7����N�����i�Aqh0#���w���!-�J�Y�2�~�c�s܌��o)q���w��%.���{�N��<
V����J��(N1�}��a�/��O�NU�#��=�6+(P�g<�qa
9iu�͙u�M������/�b��-� �� t`#��;#�%�����Qv�E�����4A��>'�����q�L$��YiN�]��$
�qun�;�L�M�ѧ*��K�*m�",��W��]����h�c��Knٰ�B����>�7�p(܇�S���t���e�T�����>(?�#��?bE��հ��:���-9� ��gJ�U�٫�#٭�����_ŋI]|���rq��wo��O��N£����\3j�ϐ+��Q����K�)5۾.+e�Z���"���8Y�74Uˠ���DP5��(I:���� 6[�60��
���qrT�S�Ii�xZ��T�	������J��P	]������}��t��zS�\M�B���d4 ���s͸/9�`$斵l��i���D��\v�i�g��ůu��_�����5�E��G{)�$e�9e�e�F��ß3;|��XA`��~+g�� Ɣ��S�L��_��ȗM_̧�Rc��/Ɯ\/���s`G�Z���*�pjr78��"�s���i��P�vc����K	2�+���N��lXڬ�ůHs�A� ��¨�$⟻����2�Q{����Wr�.	�����XlxV64EB    fa00    2110�d����_ױ	����C�
]��̓�^%�	+��<e����r���m_�ad�i��Cd
��Y7�mE�h��U=2�"$+y	#,+AE^�k9a�ǒ��Ɍ�,?�$�hЋ4J�Ψ��w!�/���3��;��"�T�K}�u�-bg13��cp4�J�x$ӜogƝ}rO<��爨f����2b[�G�˕ώ�O���`��
���P�x�c��<(zƲ�������"~�Vί��ö�j
#cg9�u<��㜘�!��Z(�.����RX��s����<7I}��a�x3�A%�&A������	�}��t�t�- "�r����O)��/c|u|iV����P(��k�n�`Z'�n�+��?v_Q����l�g�X�s
�tH�n�?�V,$�n�"��Աܐ�������KzD�O����`l`�w���F�%��h9�.�i�KDo�� cPix��`�".�kћ3�έސL��}��Pb���_S��L���|�JU�ݸ�;4H�L�t����_�e���(���m��QA���5E7-3�f���H_tު��	����`ְ�/����!]ވY�5����]p���j�P14�xy˭������.�����Ft�����]#��M��U�K�z�� ˑ�� ��j�G�ȗ���%�X�{o��@EN���!/-�z�/��!�E��64�p*وRF[��E�\Yt@3�!�i�!���f9ս3�`�~�E���M�~I_�b#-t����od���m�U�֧�[����P��+���G+
V�}��
�� 0s��V��i{��!n�P��l�6B;2�:�`.{3�F=�ϱށ&6Y4F�P�]� b(N��؀~I��>O�6�o���a�I~,%���c�U��;L�?G�G����?�p$��k5i���_�r�&��p�C��5�X��&/#yB�	��bvzM��Ҩo�wnl��u#㰆�X�Fg�|���gs�lpD�nw�,�����߰Py�:SҒ�[#��l���R���wܺ�P�<�k@�/�O}��2%�U ����y�Y�x'��蚸7���!z0�)`}�~;q`V?,A����m��Ryfc��
Ö0�U��&T�I6,�u�`v�
�F��Rm`Ѡ���=���D~�"PT���<-lR�Ρ�ܧq����i���d��2V�� �1zc��J,�'����o��K���5}p���o^���i=8P1H���)Y�b<L���d�k8(�(�)�aƊ�?Rv��B�����P۩!~9��GpQ���S���}=!1���Y��q䎅<Y����^�G�+101���]�	�=/������pMT��L�v��dY�|`�"������ZH�1�A�L��g������C|'KxF_�o� ���R^�ƍ�����7�����7���.����k*��
=^3�=���Rz�vf�J腖��mX����)�8��m�8N*L)Y�e_�0e�h����̙�}~C�Uo��(U�`T++&fe�w�=�י䠙G���5K�9�Q���!U���f�w��Bc��c�<���\�lFg�7.W��2�ŸK����FW<���)t>Ή�}�F�Fם7����ڀ��\ta9|^���;sq�ߐ"~���)=>b��O��j��D������{"��E�F�M��� @*�E�F|�P�v^8)2"���:�7P#4�d��N��Q��Y���1���a��ep��-~��@��D�l���3��#O��y�5�!!(������-���b�۵=�P<,H� ���i�w�߄6`7"�9�)=�����\�\,���C�H���~v%��	t��d���.��3�����ST�-�η��\�F7�`S#p��M5�Ъr��60�)�Q-�27pոy�jR�� �Wh��rQ-�^�����w+��@r�\�\���Q30[�k���ZS�@]/����$�4T���*��;���U#?���������X���]�x�>O:K\r����	z3�|�NbI�Cz\�h�XD(�6�g�`a��Q(ԓp��6�4��X��3�SM[��1P(�c�R��[cuyå*���lB�l���9�gn|:�zB�K�هT#3��*3@�[Oep5��]�r'y�3U��L�s�;�u�K��	x������8c��L% ���F�O"L(��h��ш��W4-*���lR���-[�r��0��a�YG��羾��U�s×t!<U�ғZu
2<W�]��T]vL�x�`l}6W�/��3g�뻬�-�fi���L�}!�`y���~;z�pM�C&���4��yf�HT���ӻ���.(��/'�!�B���ģ�7�?:Zf�U��X��)=��M�<���,oI����/�[N���CK<�$������cq�ln��m�7��5m
9?�ݬT�Ⴍ�ܧ�~+���&�{myF.9%��pQ��pn��-��RHC�U1���m�N��9�1���#HN��ڏ���}���f@�/p
;]���m�C4^��6T�V�#z�ҎuX��(������g�P�`�xs��]�����<]L�����eQ�5�з�R&�i}B��Uh��.pt���A�
|�譿��|��W:��?F�-�Sz[OXS�Gs�; �Ѓ���c43lX��(�C;:e𒬽��c8�B�\�td~RjS��N��v�so����{0{�o�ov��!v����� r4�zyz�T�!c+��%9ߤ�5(�0ۭ�
���_�n�1�V����q�����Ҽ�˶av�e�轤>�?����h�»�����>k�־0�	�e,�r����Q�R�>T��84�����(���F��t^��zր��1���!q\ۡj�?��_ńڲ��T��"���ʒ�;��� ��P�Hÿ>i3�tuG3��򉮇m`����˱HH`�~���#��/��P�qW�5@�N%����V�Yh1��G#�B���~q�>5t�ڄ���XM�p��$ސ~ٹ,�`�#��h�2\�f��C�� �m���Ǣ�4��/���e���$0�2�G���
�.�q?����/a����,��F!1����z}5S�7��`$˓p��-("PTfZ��[�ڂ ���K@��*1z�HJ|��|��:��j�0z#f���w鉆��r�9M�d��ڟ2C]��=�{�Q�J��!6��nP�08��m��xv��Z�vi���P��IâZ��,]^aO��$�ί����z�"��'c��m��1�^ꝍi%vYl;4o���ye8� ��W{��*���x�6��7���S"s�g�K�̚ᤊ �O� y�O��a��Ĉ��Ȓ\��)ǀh'Fb�P���"�����I�Y���P���n19�Y>�c�7P|�� f�gp��	0:9���u-4`F�����5����b~�?E�0[����kcs��� �M�s�Z�X��=�c��א�mu�1�������	$���$iծ%'K +��i� 4���X�ee�kv�4�D3��I�%�-O�눃h�zx	�w��r�U���������$�靵�`��(�{�P�����0�y� ��|f�Fǻz#ָvv2�%r��3}G=��pFp$=Tϑ�Z�l��%��&��m4�ߚ`��fFh����x��4lQ�N��J��d�>�ܿ>(�i�=�_sĽ�p�-���$R���d��yE45���Q�40D��@.%̷vS�� ��V|j:6�Y�:P��-�8��W4�,���(������N1��:�y0ŀMU�\���ro�^���'U�]�,N�VZ�\�DS�/���a���I��ʇN��(
.jĐ��d#"QR~�[1�@��\��%���$����1���6}76}�nys��ɢ��Km�V�NFRqʰ���\��hl���.+sX�t?�����U���dtEF�(�6�s5����V���M��}��)��f�.�\�ylV6�����
���<N����̭����:�L} �UC!�~.��#5������u*K7;�%�o0�o�����_�m��L�џ�s:U��K��~����PS�=g�����O@;����b��r?/�oG�u:��k.J��T����X���mt}������7v��g1r9?mV#Gv��udhrJ�������c�j#�ӈ�����K�~�27��w�ꉷ�S�IA�r-�$�AFx��p#M�:-�z����f�������븫�bG���O�N�4qm�����4H}JQO�/���$�͈�Qx�9{K�ڏ���ljj���
��4? "�����\��:��V��p�K�����U�z���A������j���|����PE��0��wV�ZdE<N헪w~�)L*ȼ�,�����A�����ywk��.´�V�v�a�n���;��K(�*��Z����^61���ۄߍ��I�7�;Y�"C���.\iJI4���ɥ�O�w�Ϯ�9�i��p�Y�Kq����@�tz�`��64s�|���
E����N~#� ��R�`�?J������{l1��,zLYkA-�}!��"��{m���:>]�A�w��=K���}qJ�a��
�X짪��5�!SM���<��ߺ�Q���]�2KB|~�ܳ��Jov��$�`�!�0�A>�r���������Oϣ�:�aGs��%�#�NM7��S!�����^��u�mH$z[�b�h����.�a[�@���[;�P�陲I�u�U)г���|@���<�ݯ�q�h��];X(�2\n��Wm���J���(/6mh��*Ϲ�5ܶb�כNv՚0�D���@���Rʠ5�n�  O������Q��	8ma�J��7��QKi��Z\��N�`��9�-"�p�j���'��ӝW(���o$� $Q_�w-d������F�IXP�j-r��N�D��K)4��+�_�ƻи�3�y�Y����$�j��*���7,'��c o��"d���y2�	���;�Y���;�L�g�T��\�Z����f0�����N��P&(1����&�ֆV6�\9h�5V��U	�'^�Y7�������րn���	0P����op�I/��0�Y�H��@��/���$3.h�j�h-j����`�{%LϤb+�;6,��w�P�V@<OE�J��h~�o�n�CژL������6�/7Y'4^��:�� p/&��Z'�r�"=֫��y�fBv������0��z��i�8�!}�q�{@á�JGߍ���BϬ�
;� ��pK����ty� M���D�9�<=߷��
���r�1r�䊎P�#/�Ya7 *�`X��<'�0�J#� {��iR�p����WF* �d��W �Z�^t.W�>��  W���űӾ��.�V����|�@�YD��$6N��0<{��|m���iq)B,�\܏���?�̪6�Q�B8�ڼ+F�%�p�l�d�GqS��ps+��ji�4�"jn!i��Y-�;�?.9	z�"�K�Vm̀W�If�~?�)o��Â r+@�C�e<"�����`���N�������M}��-�!��Z+6m��;��j�y�.ߌ>���q/s8�>sC�m��X������v��_,�C�T�~W�u��Sѝ��+x�S���f=^�
�A�⨲��E�w���TD�l/�$�j��SZ��K���p�����q�ٷ��K���Lr�Й��֨B��Gy�ZX�����R��P���\�%����b
`n�E�>�;7�#+����{�T�=�)x��D7ƌӟ��wJ�Bǅj=d�[}R�	�6���Hg � ^���Lp̦_�VG9���d�|[8���Y/����(;���8�ge�0]LC$Y�z?��j��\b����uz���/^^�O|�-l�t�I�B~{_k�OSd�2 ����B4�Q�!"aE�(BJ��P4�I��[%�?�$���V,(�2�I
ix�?��.98�n�?q�x��,�H�.Ƴ�No��`J�!��
C�"H��!xݷ����Ǣ"8͡WM��R�kk�w`y ��:%KT	�k�:��j5е:2Z�!��Xh���Y��B��6rC�d]�WtW�7i��"�2%����{���J��՞q��)W�Q����Ka*[�y�	�wnz��ȓ�J�Ov6[�����yL�b�H���s~`bC��b��%�%�NPL�wC�*��]�:��/�Pq��i���|aki���<��T����~�����<��]��Y6U]��e��CEw&�^��[�|�	x�5���g�+�ck�J�`�ТΓ{I�Ak��{�/Y(�P種%b�*��ǘ�oP��X0�
+�?���0O5=-��J�Mdeu,�!�8L�é�q�V���aaa�?�w���Ց�U�O�_�KPfxc�4Ђ��f�*�j�W�T��:T�v���untu.�0�P/�y�ɥZ��RZ	Ψ���c��;ԉOv�8ga�!m��NUl�`��b�����j�6��6��MI��U�5y�����,:/�~�d�]e�8L��Gk@\��X��H-��dC]]�S�cs�Mn��R�]�����1�b�<5�1�:Y[d���d3y�ٖ���r��l��.o���G����J�=�Ɯ�p�)�[�L:�S�{����A�faޣ��@��]� ��u�o	�2��o�� �wm� 7~[G߈��E�M�#�%�\y՘���/�?� A�}��]���j	FC�֬ة�a���6��5�[�՞��}6)�����w-,�=f�4����|Du{O��W�vHb)�ޢ�$�#� ���%k1^Y1��{�'��������q:bNCl'v�\Z���,���ύ����2Lݚd!͖�,s欩z�E�Qm�+�5 ���˧�E-g72e���x�S��6���q����G���f���>���a��0Ԝ1���A���w�;���2P�?�m�W^ ��|_# :�&�T�#�E �%N�3���׸N�~�o��˝~g�X]c�`}Q&�"֏�М����+������.��8�l�~V΄QB���r:�UX���$�֟�����}�����.z����$�ʒ1�La����p��T`�c6����KT�<�����ӽ�M<و(s�l�~��<yD{���7�'��P���]XW�G�B+�K��6�%�<:NW%wĦq���"���jY��D�I�CjqH!��e�a�t��B�Z3�t�0�N^2�Ӡ�� Қ?�B�8�����.��F݅bx�F�/���x��C�*j~��6c.�b��@������(t�]��W�M�f\���rx HqBV]i���{+���ִ�����|����X�.J����*(G�FT�~�65��F��H�]�s]��:k �� �,a����y���U|�a,N��B��
���.M-\ܡ��.�.(UM������e�4OEr��@V�%~\�� �t����5�8<O�M+�(g�`�I(GD����7�z�5O����]awM�n�s$+i���/�"j�V��b;_A/a�@cd.4���1�v�kf�|�����N���m�/7 �vU�=��K�u_�� �xL����6m#�k��%�P�-F�j��R��`z�5�g<�q
���P�'�{�����������r���2Q=e)9.%>��r��հ{����㳦�H{���zs�]����������򣟜=��\D
`�I/���W�	̢�a�nY�]ǈ�0�	�\�B:s��;�ڳ;h��UX�o�y����#�6��|��Tݨ�GEzNR�X����
�0� �8y�<���A�\� �����q ��l���vcs�]4��9Y�ɿ1�γ��3�n������(^^�2C�z�c=��$
�uG�pU�z��:����8��D�4�Z�0��c�+|�D���l-���t�Z�g����n���g�;at�zػP� w��1�x��D�J^c�,A�ah�k�ܟ��ǐ��q�u���=�0��l��b,�f<�a=�����Xe�3�]�����y����̥�Ց��!�T���
Mb�^��J-0��Ɛ�N\����-BȠ><�j ��._Q�o� D?E�F	��$���U���j�~�q=��Pל5�ZN�����|���D�����=� ߸��8������[8|9a~��|m�(]�MÄ�������n���~��
~;�_QF�tI�f�*~b%����� /؞� ���l����! *�y�&��ā�6�2�-$E.Q�|	_rh��B�Q��Z֦ܮ1|3]?XlxV64EB    fa00    25e0{����f��(bI���mE]/	_b8F}�`�=�E �U�i���/?��$D��&_�4�B��ӛ���C=3\��!��ʍ�ž�����7�&ǟ�ߒk�5
��AT�>q��!�؛az���q�_�b8ϖkpJ�"�vu�J����=)��E�M� ��{W�~�ӑ�Qu��J��}Y��B�"?z��M�wP�#�BwQ`C���ѷ�}�v�������F	��-,ب����u,�	P�t���C��$�a'�����Ή�:Fu<I,SH�uy@`��yP>)��J�Q�&�2k�<ϕS�zA�\��.�A#��)�������P�/��?�V�#���g|C��g�4��k���	Nl94�'���6����8`<6����\�!�ؠQ��ʇ�5<����We�^h2MM���뭘�0����}����<��A�)t϶��Y�='����6�>a�c����,���Ѝ�|	�O�"b%��X��W���}���>�H^����v���5k{�yD�ض�K�eL"�$[��9�o>�����~w�.r�Ntٻ�^G��V�~���Ci���Z<���r�ʧ�A��� ���]�0�!�k0-���ד�\�ʿ�}B�R��q� c7�^�����|�Dq���e�>1����p����󗆙��!޹���y����1��)�/+5���e���h�}Z��\�	�����|��!lH����2"�!n���6�blE��^T{t3�C�C�\�i�h�>j6���R����;�lZW�$��M��#*�@���;���@��g���Lc�Nb#��a� 	z#��2Uh,��8α���T�������y>D_���$�@�|�){aK������(�&�7�����㙯Es��a"E`S��)pk4_ڕ=���|{��_���@ 6Hҹ��O��K0D��A^�~��׫H �J��b�]����ЂiuLڠ�<�<f+I+ʟL��7�����O�DŮ&p��=��ՠ��7��!��RR횅ӛ��tC��A�J7D9X���7ČZ�]�s�{���-��>0�4�����P��s6s��Fr��~N�v��:(Q9�?qE'�&Z����/�X��t���r���0�a��6�ojv�	�X�$�+Q=�k���J{żŲ?�x�p�?�QQ�4]���|H��M�������"�X]$�o���s21�]��i�,B���%�f/(ê�䅌����l�Pl�i�H�-�Y���?��U�B=�5۶80���:�B��SSߧ IJX<�|��ަ-M�V%匠��9����e���Kz0��;9L��I�V�"�]��50*4�C=������N�s� I	>IWzD�n�.���j�����ّ�!ND6�o!�n�j$�$LF��4��P�t�L������4�#����<,�*,@m��V��ԁ
`��-�n"Z@��fcD�4_�0������8Ƭ�z)���D̂�+���c�s�v��?An�r�c'*���q�Jz%1��Q�ћ����
y�(ھͷ�nz3��zU�;�4Ո�C?�'*tD�� 9C�7N'�|�L|t�_}�U��TOR��u�����z����Ea��̺�*�����{%KU\����B����'��W��!���m}��7â��>��
�H��ُ�@�b�o�7�5�?��mI��©?�k'����Z���e�9k�k�/Kns�<O������y-B_��c\+��eo�l��� T�t�>���W�t�>ZL!�T��g���f�.�j��)
+����c��0#�kq��F�`���w��	-Z*5�@+�(�r�ZI�Q'ر�4"��}ʓZ�����b�X���f��W�NT>;��C�)V����`��F�&g6�8��*9!���]3G�V��|3�x$�`5 l˶}�#$&�*e��7���eaKinP��Fi�:e���ަ@�ƞ�a�p��x�f]̕�[W����$�u����ђ�:��S���dt!�N���Xcm��)���F��#���5��\�z�D����ioJ���|L�Q�ujV�I����T��Xcu1��.�rA��$kI����<�~��~t����=9�=L�;Ub ���>4�c@��W��*���F̢"\O���4��M���ýOBM���5C���(�� B�0�:&��pZ�1�G�� k�\�q ~m�}����h��\�+�D���x�Pz�K�0���ywZ��O��ψ��
�/��Đ.��o\�BKz�A��cdu�U�)�tl�]��0�QW3�O����@-.��/g�󩵮*!Ndl{mZg$}��A��s���R�x��TSڑ��-4�U��=�N���|�%:�=4<��`wy�(�����"�z��������^�#K��14"��X-㏣V�E�ˑZ���hki;�A@��]+�5Xvr�-���8�e�[=w�Z��@Gү��OK� =3��
�~CV R�ׁr�t�Ѫ���8��P�T�`��IvJ�E��'�f!;�/p���*}���}�������b0%���a|э�Ry4���5�MQ�l���"�fW�r��
�gI ��F���g?|_qkZ}W9>w �	�k�<V�d��� �����~��� qٟ2b=Z�(1�>H<��c,����-������q!;���7P��d��Pt�i���� ����Z�}D�?�)_0��C1����y����	��B����dR�����lM4ZC^���M��eo��O)if��(�l�hh7ЅQIu�@��,#��� ��?��"�� ��<�G�h6<Hb'�p`c(|G�e0�A���E19s��F7�}.J�lPG����<�y�l�,���	�1�)��P�h����[<�Tm�������=����8��Ȱv������fC���D\�v��!^�Z�!+%�p��(�k��I���w���ݽ�s�\�cᴲ��&I*d�U���d�Э��X�����Q�k�skL���P 
N�_]��D ��X�UY�*�?	P"3�z�������D^��t��S��Bݏ��/�;�P������~�Ώ_~�Dt>�{�F�3K4�Yi��r!K�m�z%�W�ܪ���������G�Boގk��j��iӡh��	��s[/p����ڷƗ)J�*hō�NZ��mZkgZ��lr���Xs+��$����E��2�ܠϨDO� K��h�-��FAk�j�|����V�'�a��e���������1T��4]�����X-�h��_��U��4@p���~kМ���\rES@�o���r'iM�`�2�z�-s�_�e-"��f�:2_�$_���~b:C���|�Vm% ��������.�8e)�p��FLB��l�0K������,����&o-��<qAvg头6����X?e���}o��7rւjz��8�?C�9�qY�ZsG��@��PBv���Oe
m11f�	�5yer_�J�Xرx�(4lJQ	�eR�K~������t�!/n�V�U4YV�@�#d�􌰁g�zkkꝐ4��CG�L	��ւ�j�ѵ�@��=�fRI1�p�q|o�8�]O�HV|exar���+�	ИI0�N���#�>^��o0W�O3���=��ސ@��Nu����/];�My��'u�WOM��`ō=�|�\L��LOkhL1
�hs��el�����o�$*D	���s;�+�4>V'�#�'����'JX��O�Lb����E�X����(<;��.{��:�c���I����D6-6OЈ��1^j';~��Zh����L2�g:*e�+rۓ��l?T������������Ўڈ����uZ���qq�/�E�\���%�9��B9C�X4Zϣ�km@���a=Lo	趎�2���^��o+�5�
D���~�<g�Eou�1���_A��*����lK(M��T��?�;���r��S�7���u��/Q�	��h���ST	P�^��9��n��YG8�u�%'�>�Kȸ��Yt���.�1�#�վ3p�6;*|j%ts�14��;����׵1������3f���a=|��$A\���V�����1u�4E49{{���u���ܚ�ߵm�h�W
��@�=�����)p��|�?æ����~蟠�#�O��g�(Ҵda�3 �R�V��)u�~sr_監��N��۶��&H#��~y#u����Z�.kؠv�b�떾�p姈��O���Jl<�ra��t�1݁�	�~�Cn,�}��#�X;֤m�4��  ?�y�)���"�l��N��WS��]����)G��d������ӭ�����|������zj�ʇ��ϳ�瀧��w�( ���6e�Y����b!���?���:�B�#���m��w��l }���ΰ��LQ/��%��>�`
������h��ڋ�dw�.�`��8ț�@�R��:3���?aAd�]E%�q����U,���������*�;����ڋY�HPXQ�23m�oOr߶�i�(q4�*玲�4^���֢�w&�L�wN��7Ò4EZ�/��n�F��ZBb��،�a;!$�n+�cn`�L`�_�TZ�u�{���>�.����h|��h�&m_&���;7�qȱ`���t�1"9�|%�����sU�����S���5��A�Ȁ��'�DƩ=�\;aH��X�'���$�!�����U�}����y�\Jfk�z��jp�UFM�!��@��G$�y��כ6:G�[_#F�qC[�����)�d|����U�n�^�eWƒ�N��L5�����2��V��:V�t�P����9;���^�Я#�ڹ�*�굶C!^��K-��xP�hl;�D/8��o� u�LMU��Q%A����wP��f�L�O�=����)/Ē�[1����
+�����5���"2��"�Fm�S�1���_P���P�TJ_ċ�tW�L,5��7br��wH�̏G��B�����O�?a������j���7U	/ơ����B��l�Uд�����zۡR"(HoG;�.��!��J���nC�IрW�&�b��n�'�F����o�D-P�e�����ҽU+��C���F����os�>�D�r���7hd-3��{��ߧ�c�"�7�b����7u_�_O�޻ϖ[�`��Mj�5"X�� ���:z�䓿Ґ�Q�405r#�T�㑩�8��B��d�߻��XnR8��� i�d�u'�߶�Q�ɯӁK����y��[���Oӽ�3^��3jv}H�ѧ��a��Ffr��S(O13t%�٫<(��d�	�H޶���"@O�ͰDU��q��@��-_�?���!Td�[Q$(3%��t��}�A��^��B�*����B�D҆.ld<��^�?�*���E�f�;�O˧� �8F[�GS��A_�l*���ƕN�<fA�\���B�l�ޟC��M��7���m���Q,��Q�R�qi�s���WNO��8�^��U��]?�:k����P�R�7$D��v�ߦ��tU.=<<��p`f�2�敝S�9��鑷iD�(?i�q�Ԇ�GoZ	F�;+ �v|~��ί�h�i������-V]�q�dZC��$�m��q�t��&NVyud��ȼ��oHޟB�ILeV�$�V��iom�@L�ֱs�>�dR!`B�iX��a�ŐA���.���H��srLi�]h��UjϞj��`.밾���=P�����5i�$�j�G��<�A�!ݟ�;��i �5�saa�����Y� �T�s,>�	���䎕�	"F{¡ku����&��߆�ޡ2U��t�Q.ݕ�ܬN���A�J��(*]sr����r�����p�%�\^��?a�O���~*;�˿�6�:�̵`솁�`��c0���X�0�d�>:[� u�+�H�$qzB�����|cb�E�}��Jx�l �c��[0�΁��*t��H��{}����[�
�0�>4j�G\�J�R;J��]~���+1(�>o�h�U&�������#B�U�j�I�?)b�b�}�:LץNlyp�MKX��ǿ�:� �A��r�g_2Æ�!��tb�a�u��Ъ���\�EA�A�
�$֬��C�K�R�"�m��N��k�h�=���A<��ԇG��R5���놧`L�ׂ3N�LF��ױօ�a�܌�}�9�b�Z��/��a����k� �4_.Y;�
/(�6w�����IQT�"�6a�#���xB-���+��}�詖�drtL9g���	j�����  �X�����OK/��"��'aJst]-��;[���z@ �?d�^�������T����Oxl�ʯ�i���V!.�����R��]���9� 7c����u�Y�H���X+�]�dm̬U�^�6|�[G0&�,Jt�n��Z�l�$��ڵS�&�!0F'�[3�/��wy6=Jˡ����1�>=�m��=���vU���A
�.�����:�kj�����9�	j�)n�����Ru����R�c�lz�~��.ٶ�F�Ζ����\�-r�c��=�n��f6�#a��dA����y�o�;7�����H�q9����EkhZ�Um�g�7ā|�`���#�����=�L>,u*EF�r8�� �B��D\�Nq@�������E�?�32�l�w���L��.P�-�4j�](j'�3$�����R��{̆R���UX���4��B� ���+U�~���DO��No��
#�B�y�<w\��q��*��j��<��6�鈮�S�}�{��7��BP�3L�GD�\��#k= �����>
ќ'؝l�iWSam\s�MRg|��-f���a�쾖N:Z^�W艖�!�sˍ��k��l�Vx?F�i�����%��d#Zx����+�����Qft��.I�O�Vԯ�1!�o����󫧍ш�p���G����c��0>v�3�H���fV���u*ц>'B�PbZ��.�{�勃�-9"e�<��(�ިBX�:��͓���>o�蹾��h�];
S�T,0��Q;�	_���"l���j p��7b}��	�6tjk�Q'R;J�?_��{+Ħ�o���c��"s(�1 x��KD9c�޷ ���W'ycɄ2!��IDr$6߯��p9�.H�kz͵R�8�j��n��s@c�-Cg�KԿ��]�J��q9�>ż>XW�Y4��D"8fs5T,�ޤ����[oJ0w���*�2�KQ��a�Fڹ]<8�� �W��u�������)f�۷�5i���o4 �> ����Å�/�*i�ħ?��������p�ռ'J�/�V:���;��S4X�E.��[������z.$��Fⱍ�UX� v�{�a��8�� )ۄgX�/uނ����;i:�t����@D��g*�X�[���!5[��������23�ข���G0]1�W��c�L������T^���c�}��w�-)��tw]u��X�$f�њqV��R(�^���u޳x���|ٯ�����+G4RQ�+R�ήN��aYԇ*�r���S/�q�����M�$�#��ϳ�Q�|� ��L/������}M
��!�f�;W�����E賨~	��a�,ź�4����`�E�(ֆ`��'yM \������y�'ćs�oB�U�!�k=#�-s��[��X��[�`���?5J�-O�����ߧ�����kB:����'��#���a���`t$
G�YVs�Ӂ����y�&uD�X��q�Y�/�­�w�Y��+7c���<�R�wpk���o���7X�ԕ�\��z��3�E!�g�P}�>j�1�bi�he-��c�m��jK��]70�b�GK�y�Cz~�I������P�q7G��V�q��~0Z9�:�o*%(lFuy��`f疞��L��������{����BN}�zu�������
����P
�E.��(���
�j�ϯ�1�:�I������А�a�&F�֋������,���R5*���# �u��r���̥ʶ�X�	l(��b�x�3A�����%2!+��Ȱ2�R�5���������&������I$�m3�.���$�rk�4b�-L����!e�Iq�B������bt)�<(zc���x��Ĝ��F���*�������i�vqf[��t^Mی|b�k┦�Z��s}��v��I�� �n��-=8�	_���ah�� �bA�18�B�B���K�%����3���e_=�&�B�mr�7�se���aZ��-��͹���wzj����ץ $�n'1�?��FY�L�'~%l�v�f���pv� �T�(��b���J8 ��֨��+�F��O�Et2����u��3WX��cp���S����N܆�&�ϐ�3���NN�aos�"}7H��\϶}6��?G���� U���p��U>�}d���q�rF�`��Uo,E/c���=YK����U_h�ҁU7Gn���Dƹ��kh�:��n4��9�r6���g\��@.T�٦:h�s���(i��B)��:*��m	9��\�B)��6"���$�G�r?���_zA��&���g��܄H'�`�?� �Ӿ�N�J��C�X�V&Y�0AXZ'1��_�_CMXz�P��h�����G�)��>�U��_u�(��tگ���ssjb�9��A�	� P�g���K�ߍp������#����$΢�4�5����,Pt�#ӕ"L����q�� g�.=.E�j�:Nڙ�����
�U�O���'�(d�F�c,:R<~
�!=!�` �E��@�݌p�����ݥ61�)q�nf�v:����^iF��r�4�~� g���g�Y��L��>l� ��pe=��c��V���=!F`!;�\Tp����u�)���^R ��miǠv��]SyiֶdR����*��E���e)�t0��}ʫ�4���򎏒��+X�u7qS�*��Mb��KG�J/7�pj.�m�T���L�q���m�Z�s��o-�>��%W:w�Ϊ��}<��?���b�<����a�~��� C�2�J7<��+�b�t�����x5���x�����L7��X%��`3+�n:�t�!AyhxW�&�FqZ�fB�Z�lo�h8-�5B]�/���Du�H�������I�E�{ʼń�蝢-*J�/�7_�¦" ��b��'��P���$&7��(*���v*�\i���UHpM @���_i���<"ֱ�IM(��G��W��	B̈־���b��4�6Z#�� T��t8��_i���?-+�ԋ�W��@�»G$�K���]�"��Ж�G�	=��>z/�+kj�;��:�*��|��Qۡ�qK�:L�F��"���c8�o�PN
bR/�t�O��
2u�/G�P�p���t�و ?c䨓x{�+鱵���>~�E�����Í;�4�N��jfMi�9�yG����n�7�aZX��^I��`�BϽ����XlxV64EB    fa00    2440�Kn��NӶA�29���nU�[����Ϯ���>���{j 
�������K��~KY+��ΰ�Z�,s�K��,ï+i H�)
N1*!C_���ZB�4D�-�1�7�Us1s���O����D�r�p�Q�7�M�o��7^qT	g�UN
 huq�����-U7|}��8eXz�˦��*ڤ2�o�/G�҂)��7#�Ws�8�͊���1��	RFR�)�ӕ��B����$�=�'�c�Z$�6 ��Fҋ>�|��P����i��Vm*ϼw[֩]���U�<j�h��� eq��Y�}�jv�@ϒ���RV�J6���)#]F;�U���%7e�q<	 �P���[�/f[�-��ҋ�D��e!���0��j�C)c5��ȰOC#ϩ�;�~s�FR�f�#�\<v��n�ܩ|���g������sqX���/�J���ݤ��,MQ��!T�PҘ'���K�D[�`�.��6�Q��/|mW��Zd�ܜk�[`�?�� ]@\I8'���a���&*�1N��)bP�u@��Q��ȵ|]�UV����/���b�����&q?$2���k�ɚ�m�}{p7H�e�|!-���]�vcI���c��(����߳��KKi'.�N�1[Wj��oˠ�t��q�
�6�����!!f��8��w�E��⎏�P`ើi��fw�v�r�C����~3�[УoʅB ����6�]�s5�m�Պ|k��`�i�$#(i˔{I��~����A�t
O��3Φ��2����ʈ�a�sɭ����6�[ �������u�ҵn������`�$���.�(#�8٧S�%�yu��|��\����}�Օ
�)���=:E��;[|��}���gP��ZY�U�c3�I��#��4�G��KD<����h*��PN�[�MQ��=�@u�ͷ�H��q�(���� +�%�f�#���+mÄ֟��o~��E��h�=�ji�kd4�)�ÿ2L�Qi���
�֓����xJ�%İ�D��x�r������Fh��G�H�"1��)��*'1����1�m�ƹ������BeF���`��uP��{��	 �_�������Y�~y�SCRS�2�K{G��,Ӹx��ԗ��e�'��a֝3��(,�z��c�(��[`�a��W��@��+6`kvIa�B�,қp� /֪Q*.��"���b�P��a�R�V��y�3;Z�|�R���Ia1(f�r*��)��A3�Q�5�2��,�`����.�7��Q:v)L�\�/Ĕ�ي��w���l?�ɓ��{PR�Zn6`%�7���¶|�Ye��-9�����(���������[���	�	����K��T&"욱A	q�F�'��T)�S���u���?�[�mR�ո�����:�+@���oK�2�ೝ1,�x������6��ó�}�|6�,�u~G�U"ŕLU��̋�Ր���"�m�ZiՒ�y�U�����)$F��<��p�-O�V�F�׿����o�n�8v�R��k� >�o㣝����tr&�g�4B�)�#�ײ�Hf.��q����j��0������ ���P�{�:�T�\8�8���"��E�6��$k@�Ws}��}�|=:'�~��c�>����n��(@�R��>��!�
A/���#W�'ie�L�bO H���#�xJ�煝K~��.�;j-t8����=:��y$s�e^t)��?Hc��lhD�d-�Ǚ�� ڹ�D��6�-Y�Pwз�
�stYv��zP��f�;|�`J���^ƾ:��#�[,�=N�I������9�a���w?֢gD�|���B�RP}6�4���;��/�+\�6�GtP9G[� t�V���De!m=C��R��B �B�o�<_mFfv	�9e:��h��>�P��n���S:�&�'UH��(NYņ��nb�� Υc�dЗ���yHx@i;U������$���kC���z�7���6�]�)�9����|6�<)�`��j��y��PG7�9�t�4(��Y8'�#�8�H�F�%W�э�R,�~���`�������� ��-3��̍U���H,���NJ�߼���򔷮 �����Q�/ɥ`�V���і���f�~�cH�%���+P]W���N��Z�4B�bI�({��A�8.o�����qeYmD��8;ږE�Hh����G���Q��tl�������v�l:��O_�b?�[�$�X5��'��T�k�{���)��9t�ю�������o@b�����f��pTF�4R���%!�bؗ�RN�E���qH��휶�	�R:��t����H��0#����u�yk����6Ƞj��Z酁��0ڦ=����I��\���F2��^Kg���RK�iF����@��ު���{a'����h8 ����1+����!Z"��Ȅ�o6����n�~S9��ŦQ}�����?f�H�9�/�5U��Z�E"**��h� Ɐ�a8�]-���:��*��l�8NC��u>��枫�q�x�p�y�:��2|V9~>�*:�O�|̾�~|߻�!#̣�b>?mw�|�zr=0�R���Sz) �Y��4b�b����_P`Bg������� ��V?�_1pf�ţ�C�;�^V�Qp�W8�ı��Wi���Xb�vp�9���[�O��9b�w`[ntCU�Z�\�� j�<�Bd.4�J���ɖM��^�����j&igxՑ��]�O� ��m��?]5��~�ݳ7GÌ�j��f[1�DϺa.��6_;鲼��.�jF] vu���l�>>��~s�Ez�ǃ7~3���/J[5j�+X�����ubE-�d�
�������	�و���PS/O�`�'��g�dO{�T��Ң�q����A��z���0E]D��K�H���R��%f_༘ۮ׎Bl���+��!�H�H�.��ĩvN`*s��p]X�z��|6U���5ۨ��Y��D(�9���0���`�Zf��.����y��!����������5ơ<0�N�1�"�(osk�A��Y������m�0�kg�-q���/oqKT_H	at�S΁��MT�k}5T�u	]��;w��!f]��-������N2�\���aZ9~��IFA�}�N?6�f�*���Bi����j������˾:FV�8�(�SIV����P+[2�g�y�&NN)!Mz]M��]<�3�:��>��=��p/n� �U�8�������u��I8(����X�aE���n�H����[��8�n���R�
�-<�[Gǯal�V�+��9��Gq<��~/@T��?�Wb�,���^&
�n�#nM$�y�;�2Y��n�����`-�;�����4��Y��H�J����I��u��A�עū)�j�������~�����_6��2�_��]L� ��qZcʹ��U ��AG� 4K�}�،\˛A��7�f�C�h���/�p���	�K�%��Iň�ix�ac��;W�cK�G�@}`�u��⒰7�12����̧��Ȃ�z�Sz�]Ld/
9���z�щ���,��$6�Bꈪ�"�}>��~�y�0��P�_��I�o&�~k�F�8�ʴ%6�e�
�90���K�p��0���GK:���W~�h�㲦hN[��kJ�Y]�]+���įr���;^�z�4��~�Ș�*a�9���]�X��Ϗ��ʺ�-m������Uu ���|e;��P?cv[�#p�f�?��$w̌%W�t�*��ʒ��_���i���ye?l��|����]�6(r��ǋ���f�+��&.�!�,b{q�@1KUEF�������CfB�8{1�����\���Dk7�r�"��2�%��)���{�4F���cW���Ak�)mWe�+�V�����e�|�DHyv�Xc�Zx�뻥��q��)�\�:��&Z#�B�����b�+�%�\BTw2Y�	8�j�+�;y�5�P��Uh:�-�CH���m&���L sW>Wh�BBy��4�z�/�M�&>�?�:��Ѥ# ����\eދ�(�Ԋ��
���gT?pb��Y;�،��r@��0�d�.�g�?�%�}�"��D�2�m;�=;V/|�F�p�67�R��>�:��Gh�M��eCm��cF�#��@+�,�y���
2�6�_��e7΍�Y5�i Ԇ��gg�4?�KB!Q�VHz/���?�#<pjp�A��4��о	`�=	KBE�N������+�$�QU��T��C_r���[�} cWZ%)0�z{�Ȅ7$/�1��{�ɲ�*��$���]V)�҆%<4��q��_�o�~��Gl#?���U&ft{�&���Lo%9�� ����?Q�$�s�®e��T����G�8���������:q�w���Ӧ&o[w&7
'1�	
0�\(�A�)�+`���h�Ks�N�X���,�ryAzͦ[:uKН���kb�
�ez�����V�x��vJo��� X]���$�bo�C��*C�W� ��Hs2/��d?�JB���� y��E�̽T�A��y>�vxf!a��<nb�^/@Dh*f�T+�R#�D?��|����-��K�ꖲ����ϐ�lЙ��4��R$t��8���w�qVy�b}��oi�&���>�� g��z��l�FI����4�q'֛ 	��C�s�/Fe�m�(�٧��t��C4�]������z0:9��:� y���J��iY%7
I��烨�i,w1!��6���w����w���mq5�oߌ~]�٪��j��)�[���P%>G���K�lh�3Tw��"8�c���x^I@N�z<]l6|�FZ����r���9p��'�zu�U[C��Gɝ�e(�g��5H�c"�h�`R/�a���S�� �]�!����b�U��N�����b<O+�1����b35�H�\M��'��1�㤯?�����Ԡ3�-��,��o<c`4�$(��j}5k[e�ך�Y�@$1���~���P����zi;g:�T�7��p�]A����5�u�Q���o�4pxB<����O�����c�{��XʈS�;��W��-X�GuMgQ8Vˌ3a�}:ҕ���h9v��Sã8��0#�MO+%�H�LӴ#��؎T�s��2��|���0dqF ��V:� �9<{��c��e��#�_˞�so��CoO2R-eW��U����uO	�8��xx���l�C�<9K{><������qn�bi"0�%�݌���C�j���^e��X���A��:��HU�*9�j��Q�������GF��z��?IA�Z���&���^1�z����Ё��>�a�	�	�Q����T��ĩ�&�j%݂����f�5\PZ=����*�"/1,�A�' �7S��d�[$(�<�)p��k��d����s ��ׇ�7��4�u����)�tbs���Es��pm�%y�Y�}��.$\�?Ur�ځep;7g��?KR��B��z#�G�Ed>���Yw�Q�k�d�{:r�����Q4������%���R�}�])��<�5�'��������p���^��YM�K*2�������$Q�k
����
l���?���B̀un���ǿ'Źp�#����c�wiO��� /�IV��L��@?�l�lv��4����l 티�'OH����!��.u.LC�$J*�-�`��p�@l4=�G�}��W�]���0��do�x~���6�X���2��������	!���_67�
�zU#Y5A�-H�]���aP^�J/^-?h��l%m��!�?D+?X S��
Z܂N���
G�j24�7�>S�򛾜k����C��¢Ƨ�ߓ�?�f��jiڲ�����  ���'����~Y��S[R�A����٫w�0�b���t�������,4�Z���J�>:�1��F�����
B	��X �^Ě^S�H��FWB��r�xk5F�CRo{�\m� �}{{�H�o�k�/�-��#=a��a_ѧ۷;3d�"h���0NqI����d�v����w~E�Gj�BA�i�5Z�h��{���$o�_�ϒ���g�o˃(�
�oLrO�m����zo���e��G	R	 �-�]�Sb�zT+���K.��#H���T�*NGA�|�a\ģ�E�=��e���q�b���������?M`��>N� n�/���"*SYt�OU���5� ��@:�]���s-�dx틩eDcr'hQ{g��"-��`�/�R���L�Ⱦ	l4Ә�4��RO���$�*!a�\��T�l��hB����HчMn����:x�T��S~�����8�Ll0����j3�SJ-w�KJ�OӜ��\�`��=�~��N��z����ކX�/c\�h�v�#1%�^�?���h���2�9��I��b+����ąy�){���l�b&��{����#���It��p��8ଐc!��_��LLѠI��Oo
���8u�\t�tYE�M]��a8�(�ܥ&���.��5*��"��1��p���t��n����m���J/�� �a5ө�.�{�M�bok�O��G2��`jt��Z��� ��;��C�❡c�m6LE?C��.����JE�Zp!BQ�]>�v]u:*�|�ɷ����)�U�ƿ'�g��o���L��C��é����)��ehmB���y!����εH�).8�E.� 6����"6�/�=�]�6g�LE?տ#���? �����>�]��>��eF^*�,dg͸�NY<߄8�(��러�����TX��冣�U�Pf,Nkg��0��)!AE�D�XC�)+�ȡC��B@x^X���� �`N�/LT=`���4M���h�߀�ZI�*:+z�� ���gDe��c*�%4���H�D.qĿ�C�%q��m�E?.����6H�!%U$����ƒ�(���tA�j4-��%��$xʨ]���i��Z>��v���f���-����� w�f9��;�`f)���pw�����>�����sv�\썮�Bc6;�h��KƕH�;I�
�|�`9���ުRru�ˮun�'�ˇ���2S�y���lL-ڌ`�wǰ9��":��	��D7$wj��؝7���ߧ-�	����M~v`qBk���%4N<�8�Lx����Cz�0�����aHН�2���	��h�pc�g��g-���G�g1|v��7b̀@�6V��}X������ҜfѢ�3#�m# c��V�����b�R	D3#����X��-cw�����{�MA�����q�УSΐ�ϊ�煪�iNGK"x Nc��=k)�uO������4l�p�Z7����m�� R�����Z[T�_����:�҅�;��m�r�$��1����o�- w��� Dc��M8:p�_����mP2��Mh��(�@J�k3^��|XX�!�ơ_�	="�"CqẒ��`�'�>�ĥ.�L��#}�2���%rt�(�<�ds�P$(14���{�V�&a�78�`����A��Ø%\�l��~�:|{�r(�8zFU�=�X�=>�rL���5�v��͌�P�����77��"�0�1Q�#�H-ʵ~B>�ⒹB����덪���p�!�P��0�_k��U#7g]�L�G�G�樲�b|��x%n�^2�A�I�Zο:�x;��-��`0ӕ�'�ð:�f�%ꖙ�4aN�+�-�nlq��y<�k��x_w8�p�s ��:�j�כ{8�r�r&n�f�q6���lҬE��cp��L����w|39bhoDf�-&��uR��-ʵ���4㟪oA�N�͘���L���ӞKT������5�k.�&�w�ϓIe�{ՇumL$1u�i�U�^W�M��Ǘ��ݢ��\h��^�?�!e�����]�w�m�>���29�*�����I��D=Z��<^�Q.b�sx7�<�I�?�N'.djQ��J]���}_��Ѩ�Hz����w�qq/�q�!�d�����7�5�t��f[�Ͳ��NȒe���hK7��1;�`Ɉn�P�="�Wn�.!�ڂ�{H��^О{���������Tk=. m�e=�/U��e�� �ţ~p<�W��}/�0�Pl�K�qU-ǜ�������aTv����3�v@~s���D��vi�I���Az�x��-B]��_{6�l�������������QO����P17�5��2�-�7�� ���_�������)=�Z?��7�y�?�L~e�p�M�ޔ�Jg�4Ӕ�U7�[P~&�;��N�A�Xm��J�|"�S��'�J�apShfA1$�ܗz�A��M�G��Q��+
!ϰ�y��7v�!��X���SA�⏝Q����N74�7֣, d�����K7�t�������Xԅ��#���sx5�.��ޏٌ��� #�V�N��ڳ]JիX�ƈ���(@�K��w? �X�w~����R��W�:��c�N޺���@�/^ɑ#���K8v��%�C.�=�--�R	HK���N���D��@��
E�	$k�#�9]��9�Aǈ� �Ӂ����	OY=�b�`�R_�e)v�ˍ�1%F���pmƫ��7�
����W�1n�{������7�������m?�m9=l9�.,��VJ���e�7L�P
$I���R�cϔ�g�ߟޯ�����<��H5c�������}!�r�EP�ҡ�ޓ�pF��n�#s8����"���v{�R����Q�o
�k����iV��+���{��)��BnоBI��bb`�>�ѣ� ��B�j�m���Р�)H��]�G��G58#,jB~�
\Ca�&_U��f�T�] � $���$��@����k�r�ͺe�ɥ����̡|��)�ˮ�Eޢ�k�#�8FL����R��;>��\ퟺ�L���GVQu�`7��b�5:��S)�hɔ�ͨ��D�hPU��P2n0�0Qc�;�q��-�BZߤ�5�����jol����=R�u\2�'-
��L9���#;�No/Bw�mv�K���"N���k��L>S�}v	~sӴ�C>�����*���8����XlxV64EB    fa00    27f0��fru���;�n��|~���}�',� "l҂X!�NbnŃ���I��*$r�e�X���'��	�{sHG�����XL��� 퍿k��u�ؔ	g$�x�4ǝu���(dlU�W��꒰SjG��r���_�!��z;}h�w߼��~2���9~��}��:2zҁ�B��\��F�G%vEr� <��P�� �� D�{�n�x���5�_K�,��NwDo�*��Z�:��f��:��ۚ��9��<j̓���w�Y�	�Lle2�oA~q�����O�߇�Le̬9���������G����;��u	< T�7 �Q�!��t�OezW���I����Q�}rN9�Xc�Z�8�p��s��"<�\}B�oy��(����л~Qj9�d�5��@r��W4q��8�<IK�K�[�����|nSM9�_QH�)�a�,`F���>0�|��@3����¨p� �hg��qM��f&�f^�̸���߮��ݳ��O%�eW�xf �V�,̉����`��9�L(|���>:LЙG�T�%��d󰓭T`r'i2���
;�S�1�[t2r+q�Uj��r�H�rw��s0x_�u������ �y)�Q���4�M�:�
`e�8� >���'-z�pa� �U�jk���H�a����{O�� �m�؄)�i� H�]��X˦�x���ng������?��l!?��j�u����`�q�~"�&��7�7��������r�O8{<8��q��;�ĕ��.D0��E�������k��sj� �2���W��T��IX*��4�Û��N�J�q��!)S݇#˗�ݪF�0�gf5���s.��
#��f�~&I|�\�wD���E��I�]�iP�%~�r@M���1.9�^k��?	1���Ҭ+�ό�Á��=�U67��!TtB{�m[F1Ba�c����̮-#��\Dc���F���^7���l!�j�"Qm&�[��|��7�$nl<�8h����ba�]y5��|�3�q�2���&��R�!�U�KR�\8D��6'b`i�0ۻ��-��<�ʐ�x�~������U.M��߯�:��dG2[��w2f�V���+AFpˈ��Dv̸�+ٯ�z��3����(�C��}j��8D����pt9Kf��!,��&�>Kgv6�/?�Bs��E���S�;��NE?����Z������]> ��E�&��z	i39~dse薃&���a���ajM�I ���s=''�O��W � ���?��֥�l�͗0!$k��E�@�C�j���t��n����Uv��2��P`d�F\���4�.E�1���.��aS� ���Z��:cx�A��T,<�z�e��}_����-T�|��%�- ݞ
[���SI��Q���+��Q�,�0 �7��K�x#d�>��m��	z�G���������WG4�`��r��{�ƞl������F�d����h�ԇ���"�r_Ǳ�Ò�B��Z�*T�$�6��� C I�i�~̠c�B/��3==� ��[��jjHM�� �-o7�|�i���c_�l�Y?� '��]Bdw�W�ȕ�p��q���jX�ޥ����Q��9�YalzoK�7K�߲^�rśa���Z,���w�Ș��s���Я��``B�R� W��X\�4�&���O�W�B�P�/n�ʱD��������=��ՠ��RK��
�K�G�@!��RB���oC�6�NX�P�!c�BF��-�G%��ϰ�=z���m5W��<���k���Q%�2��^�65��������c�23�Wp�����^B-���<�An�(M�5A!�r�ɢ�:����=횝��ٖ����rp��x��WC��w�hGg
7�T�5���
尲Y'�}3hNr2��v*m�߇hJM;/N�|��C�OŘN�5ۡt�*,���p�HaY���N�F�����(�w�u��D��Zq�Ƽ�`�8��0�]6������[�zib�=�c��JZ����o�ڸ �d֊qx.�@�}VWU
�0�����Y�7�K��`0�'.�3T	ش��K������3%bO'��H+����RカY%cR�?��e7��CeP֛���xM^49m��y��*L9NqS�����e)�5\J�:��E.��p�#I1=y\
2ï@�ϴ;~)�����|l���`ƅ�ac�a�PV�K�q$�$ЭM�6}-����@oX*�<-R��1
HOAf.t��I�dl��F�?g]��'k�<�t�q'�8��,��k����F�
�ߞ��<������$	�7��%��)G���9?֊A12ơ�О�˛�O�Ƃ�hk6�5ژn�\����s���9�u���O�
�ޅK��x���\��Dð^F�ı22��~J`��3�J?b�� I�f߮���%{]"��B1�&ԋ���Q�#�	��%D��v��v�,���all���nyw�B�\���%�߱�M�!����p�Xo�ׇȑ�����$q���7�9CA~.�dUf��Y�XqYw^'�ű��}��B��Dn݉P$��BM�* ���x���(����T���$�al���w���w�;/�h1����S�5��l�%��o-����и�PQ�eg�aC�D��:3�|�f��q�:ಁf�J$9�_;��d��a�7p����ưZ<��sd��nA�4]�܅����Kt!Ԋ����j��́$;=n�� �_&���gDMP�9Y��(����N*%du\Vκ(��[S�����(©��?���"{��â>��T�+�Q��9��VU��+�Lkz&3t�w������'���f���8�=�8b���p��O#�L�"A����8�ݬu�jx���W�(
�zW������H�r�n=k�6]�Q5@�\x�`��E��6-�b='�˽\)yNJ:����+g����SE�N�6�ۅ�Z$��ʕ�AF�O�X�C[die�O��hs��R�җ�f�UY��������8=���;L}(�h+�,�#��xq�o*� ?g�
�y���r1O�O��IE(B���鞧�pX�W�*Y�Dp�k�Y�)��sY�����UuN�
�j�)�Y(X�)z>��R��d��]�j��1�VY�֗!��A;��ZQ��fp-xt>�ש
[%	�f�P�MO�-|��9�&�:tU,��>���`qWǯ�M�GG��xD��Xj��C���DE�p����2�2���N
�'����4U�����o�U�CK����-4p r��$�ެ�C:��\2Cw��Gd�c�'pɚ@B�NQ�+��u����۫�>}*}�	؞�}qu;_�?E�$n�6��qz�P B��諳�-�>N�H�o�P6����ֲ��Y��
YT�19�߃�-������VA��B�E�5pBࢊjHA��i�ˊ8�ZX��ń;C�[�0�F�Eq<|����Y*˰�7��VQČW�O?a5��Wb�Hvs��uJ3|�e^u�E�g��;�d�vy���=�GX����le�s�JWMRM>��Qy��/����(}s��?zSp���%+.'ގ{�D�)�W(�]�F��R�"��r��KY	_j��`qo�ӷ��%J���L-<�hB�e����s�������wkn�E=$|�#�,S^�R
-���!9Ay9���Kz2D3��F�3���[ ���bnD����3SY����1�Ľl��G�m�G�9���k��Ӓ�#�k���ڤ޾<2c����Axܜ��?}��N���H���s
���ej��L��\�i1���*��\/�g��ɤS�n���7�ؠ�N�MTG�>.�y�]^D��^�N(K�s1�H��`��Я�x��ڗ��m�D	 ���(?oXC�6!S2U%��.5�;E('����M=�:�T�^D�{�E;U�g�^@��s�3z��s�~�=�XǨ)?��C8��^^#��������G���ga2M��y�r_(yi<3C�u<�`\S��#8�j㡄��(!�k��dR#�?�Y�p�t?�+�6�B$�e�UB���_j�`��y&c��o��	xP�Pk�'�N��nD���"���TӞ[��O�p�r��,�f�ك�	\�Ðv�i�k��*vG8.�ܜ�hU����M���}��v������d<}���g�a2xf!$3�8�$�s�U6����=hH�����;��������d�ݐ�64Ѩ���0%c��R\b��yJA1�>؋���W д�Y�2�f�b��V���pP�t�	�[ϒ�	���9:kL}�,��I��f)	�1��[�?�ǲ��u�c]Q�6��2B��z8�0����)�i-E��Th�(�o��>�]�80�">�p�T��ڮ~7�d@-���T�=`y'R�گ!�b�<_ٺd�hȩ%>|����i$�/�M��RL���2����kKh!,����u\FRyW��wQXp�%��zd�N����c���y�N�?x���ԫr�i�$�x��{.�T�,/��X}��f��We�A�_�i�x�7��_8$�;����ơ�m�P�L���Ij� �S�����(2x���A�3i��H�E��j[���CK��cuKYl�:*� �u<Iu��bүa@�S�\��f?x����b���rG���
���R!���~�_*'	�2�@�"�7Y�4\��(N�{�x�q��I�+��Z�����
�)�v�)�CI�.R�>�d4�Q$ô%"8��{���+7�b
_�C2�E�.�w�@A,n�"��hI.���X\)����<Z�ƎK��2cB�*Є`08���@"B� Œ#`0��w6��8P��x`m���&:�
� "���%���ַ�~�&+~����.*ݗ����r{CTɛ���.@�zC�d[�9��W����dr�%�zL���"�,�<х~�t���xZv�(��:�U�ͳ1=�� �S1�C�՚���]��m�F� $
wB��EJ��E�l��o�T̲0�mH<{Db���mga!x��m��AxΏa��8nB�K�X�v�V��U�Q�9�\��ڑ�1�ǘK�1�׫��<o�b�ӂ.U�@oe/�m*t֗9��$̋�� ó����X�����
�N�J+�KVk?�����a�/Ȱh�+'��z0�:"��\�C�7���}� ��� t	�ν���H�8Xd�O��L��kޅ�to�DFB��<�gN*,�j�(,��pɞe���H ;!/�B!��Liώ�Ʒ���&��4s`���Mx���`�
��P(�XJ���	&U����2(̬�v{?��#�d)J�o��^T�Ν�W�q�5�z�:ݪX0�xWU�<.�]��mߌ��+�s���P'#"��Z�m���0T��u�(��Bc�ܩ�|_|T���P=n|�7��3r_C4�/!I7��U��V5G�S��eΥ�Q�L����Q@&2��Z(}9��"qq�F�tD��~�^+�R�7��i��H�/ c����ˇ��&lϤu�����h�ha�Z���p�6˄̴-'K��9���`���.����[%�6C��p3=�����c
�[�v��`������Nř�<��u�j�J�U��n��$�I|VEci����.¶�J =AI�p,%��SBث�+9��6�����������h�^�ks��J��;2��#�(.�_��_�������mq��������=]q�ڞI�?�-���Q`�7F�?nn��/������s
�m���H���<&��w :�x�[)�r�'6ھ�	�Q�Z��(tB�i�^j�����`�I��Q��R;9t����u}�wH�
[�7d�(��E��'�u��ߐ�Ru��&�e�Tv0��  �r�\1T���W�U�,$��ғ����[�/�����>��@�0�)���)�M�ٿ�џ(�%mJ�\�M"��}r�B[��"u�B�]^��1�[~���Y��7i�ZC���j�s;�����lkJ�	w%Q���"㮞��q�\I1��av���Q]y�i$x{�m�r��S\�ݴ��4�+~��}����`�e��q9�?�-l�f�K_D]��-
�<(Q9ug!_l�����#�L�LT����6N,}�����`T� ����F���r�^g�k��u�)_�Σ�O���[]F�s1�������B:qz�����rBgJM�:�R������7&E<�Ћ}�DfC�"�p'E+9�<cv�boئ/�xxo=Ve�P� ���a�@�E8�v�j�H&?P=!h
x��p��f?l;��bl�K�e��A�Q.<q��N�X�
���s'�ےkE�-
�FN�q1�jV7�u�R���e��;�����n��;��I2n�:ΙT����pK&Bn��Vr���	�ޘ� ?�X��d�	���L�m�Y,�pnZī�����aLK�G��G��;s�Ώ�4	.�8ќ�c�������y!j����L�A�D�^y�<nk�d�!,�=�,����YPXY=,b��������D��Kѭ_���S�Ȉ�`qzwJ��L�v���H*x�_V�T�.�3&�kZ��=��>_�O���K'�'�]�k)�v�x�B�bA�5���iTx��)`�-��k��>�a�K��xQ��!gi��Ft�mt݆���H�.�`�K�'��	�+�c�TM���k�������@���,��c;�l�X��֍���)���[5��r�G[Mⶊ�.�k'�{��g�j�G�K���.��w�����D��įv�� � �.�h撣ݏE�,���S�C�^u/Kw��5�i�K��v�PFK��w�4
�jF^�}�fW�j�Z|�S���� �4g'3OX%��=��T2�����f�s��-K��T�_2/ۅM�NyB�ӻ��d^��'��|^7�̘~-��|u���\���0k��dR�E*��@���z�C\�`���U������@=�!�g�O�����roH]��?,�)��y�v"��q4�D@K|�R|n)�R�5�U��A��6��K�vz\�F��.+ҽ�L]5�Zm��}�u��fհ�ݽr�kĿ��7�+��V�+����P:���`�hL^<�-���wG*D+Y�=��y4D�O��ߴ-��u:?�[T�L~�'є��q*������4����q�/��^��g\k~vaG4-�o��1k�1܎�������{-���|wj<b�ذ*�ȒӘ���Dٺ`}���S�J>;e��P_1I<ǡfw�?j�~9<�g�n��s]_����b(��}�d�Gu�X���9m�G��=������Dԋ���� �� �k%ل+OVTZ��jӯ}�t��W�3�x/`���(�l��t�-<5���J5m����U�Ӥ�G������ŊN�_��'�IЙ��=�4���WS�/=u<b<|�N#8^l��X9ߴ���r��h�P,߯x<Az�������ۭ���#,�u<�E�~=`6JIh����Q]j<��Jg�ԇ� �$4��]�C��8	ː�}y�2�a���#�B��G� �1P��Et[7��G	�J���`�[߉l�ʼX����UIy��s�~x*>�k�ӣ���X\�Χ�� gשo�!	z���]Q���w ���7�)�5.��gj��Yw�A��?�X$�#����̺�`�XD罡4}N�ں��Y����c&;vX�s;�C��}5?�����b[k��2Lw�%@G5<)��\µH{���(�,�
8 ��0b�<<H�Ӷ�~-���P�mK@3乎
��T��$�7�&��'ԃg\��kZ���K�G	X)��eKGU�*x6�X�MQu(t6np�u}��)������L����V{�N~�L���y ?w3�k���!�vs'��qܹ��el{�h�-�����<�%��)̑��c��k ��0[�<�@���QXw5�� ̗��Z}��g�h�M�M�܉�Q�c�(%�����V0����@6ᔏX�#�x��?R}��S :���fǼ�n�wi3I֖��v���/��9UI�����.�9�>�����e��&�A�%����9��u[�T�H���d��ǐ��"lW�9[7�ȳ&Ǩ�s���H�኿�p��5����HgPH#}�M'2�V�������!��Yʳ 
.i�k�Q	k]�u=�U�rP���*�nT2�Ɇ}�$�a�/��$���D��؞T6ݍ�!��$���� .�?A�p��^nꃏ��̃��/�����Y����c7�Z��������yǹ%��R���}f��0m���^c���;5���L����{�ԩ�3���A
�~~U�2��p�էo.l���	�H��C�UƷ\vq;�L��P�3D��*�,Vc�ˣ�a� ��z~���F+��F�D��*@Ƥ��/����.�q�y�y��R�	��
f�c���u�����1lĺ,�*1����Fm��h�U��&GT�f�m͒	�kp�8mL�'�<[�!�ed>��ۜ� H�\�2-�W���=������p�T�7�+��#̃��t�f6N�����3�/�돖fչ�+I
�Ʉ�Z�*s	�LT�t����]�IO�����@w���Wjl�[~�H�߳��A�J��&��2Z�3*�L�M�U�Pw�?����Z�v#�\S�M_���R�8h�(��3�e��ȶ�T�g䟑�2V4�.f�C�j:����wgo)E�~Z�/���9���?^�'��yT���~$��w�:�aZ�ڥ�#k�!Z��ڑ�O�M�(O+�eE�x�H��y�GwF�*��W&\�A�\��/��({}��|z����
��R��T��UV��c�R��@��!��;S���$�1p�=�=��2LB )�,U� ��[��@��M��r('L�e��[;����Y�<(a���^[<�8[�s{h�u��!�lԿ�\��? �˨����}db�:�sp)U��Jf���1�OA*���@��=7 Tٺ@5}>��^���Um�*�f�nTox��b$,�q���b@Tp�M�ӥ�[C:�COc߻G�d&cV>ᎌ���L K�l���{:�}�x�(�N���˕l�a>���*�ܠo��h�L}5|�n�ˢX G�� �h�_�∾���vP��ܛ�{~��*"�D�ϫ7	W��=��d�"wĝ���O$E���b�捽��H$A�.��連h&pQ����G�������RXbZx虨?�1��3n��e <#� ��%���&u���=�5�{��ɺe���I\�K��H��a9���������� 5��Q1e{ote.��J�jo��j�X�/x�$����FI�A��t{�H��מ_�����S&C�7��Cu�I5k4��J~ݶ��a��7bI��`ɡ��Z�ʛ�~@�|���@R���<e�/l�����/���+�A�m��5m7�tqn��	#�*#��^p}��wT��0>aVh�w��C�����_r��0��|=�-�
G%� �Y'rY�B��x�p
���%�u+[���Z��2��%e�>�"�Z��5�C�M�J.U�ךgGin����_2�JCy�*�'J�%��ַ���H1�^���;��g1��M$6ˋ.:�<��xkɑ%�v�b�n�0���Λ|�F��S��1��%��oU%~�������P\��&mW_p�o�h���j��~}1�1�h�c��Z>�FP��"�����{�Tֆ���j��9�?��M�~VuɶYD$M�ʔ��.�r��;��i�݃^����P�ߊ���Ӌ���)��	�`֛P�E�r��#��Xl>��^	d�oZJ��3O#�t��"⨉�睮D^LFЈ.�^��Q
[�\) +��su�'���ur>�dZ�9�Z����z?Q�@�i�}��Jg�(瑩5ЅǚEx%��e�5�s�T�T���,��<�a&�n7����yc#��Ϧ�D�D�iY�ܙ�K=֛��Aӳ�����ǇCm,��o l����Z]��Q���d�Ǆ�C���̉8����:���F�
�^�d?L	pC�(����k����]�AgX��/ g������RS��XlxV64EB    fa00    2500DH�fh��$��UB1D�����1�Md⥚))q����=ǋ-:�MhA���Gͽ�To��H���$�0�G�Bb|�]�|��Y;�P��OQ<���W=����6*�0W���-�O���r�vz-�_�ӎ�b^���c#�X9|���w�x#���>>z�5�3�����C�,��Gr^P�2�-�]��'���k�{�t\�C\)�<`UvZ��[�����-��ZI���[>���2�Bϗ�Y	 �A�(���A����<%�z	P+�k�2č�m���`R!�ǈkP�:�w�4�������@9�=�rN�������`op������Y� 0}�����Dh�G��b1(��ِ<HnCP#{~��H��h� ��.���s�2}��� �|oIB��Meͻ�
'O�zFC�@lUkXP�.�K��#X>L��r�R?V��M	搅�P�I�5�&�4�k�=mn2DE�� �W�����V�bɕ�\�1�3�7˘�3k��~�+4�p����-*I�^��8<�e+��n�ׁ������)
����}��4�vi���V��ΆGnƙ{`�6S��oAc���Xqn�k��
���� �7ިL����/��nm���p�J n]т/�|����=@ı�8뺠���"��<����{���9��]�M���1�e+5�X�X��O63iܤ�T����L�OOM���<,�L�k���^�e���{u!���ܵ^�d�� ����G\j9�w쎽�Nh��e�&��HqND��(1�6�/�+l,QY�U������î���@W&��Z�'�c���AV��)��iy����P�)���Z�#��VJs����K�{�ô���$�(Ǌ��z$��782s�P,��[��-qfQk�B���g2�=[�����?j8���
9�%|�tm���{�J�ﭹ*H>)^���E�]��k�rZ	l`��LJ9Jo(X�Ի�9L���Z�S�Vn��f���y���,��/Ϋ�Ր0�*3�����{�%������W��k�$�nz���"�zu>]�E�u3�抇��:�v����k�k�NI9l
,x�UɎzyw�y�N�dʼiXJ
�9�QK�WN��B���"6n��EM#+�+�
ƌz�����5���^����*����0'V��e� � �-���=j�4�)$�D�_�?$���X&�Ʊ(,�M;�M.Q �[ȑ'{�>t)�^�w�q���P_�q�4�\t��ܗI�K�������O�iʝ)�y���?N�3D��̪�_�J��V�l-)� (X���vm�tW>���LT�Z���l��k�[���ۧ��ꔹ���1�Ʒ�����h���0a>u�"���V(hErϯ	�I��%8��[���� 8�=?� +�Ԏ��7:���,�*�n[j㮹/,Z|r����Z'{\�Ԫ�
�/�Z�g��w������K��hz��+������� �����[0�Fm�C`â��`�%�?�J"�5��X�� ?��h�ꉞ?���E2�ThaU�M���Z���o��A���z�����(=.0�� Q�vΠP�I�F�����R6A�83��j߁��^�!�zHQ-��`&_r�H���?����'R�տ�5����B��&j�*J�U�cB0F#������u�_'H�9&��7J��ݑ�q@$��UZ�KU��FU]�����{@FaM�:Xh�#<�5;�:���jjM�>n��.���6��S�������D�B��>�_x�8,O*���Z����/����1���VO����ch;^�*O�L�by?�*歺�Y��cr3��
/p��}������8�m�l�a�H�iWaƎb��۳0ҹzmx�HE��"��S���Z`!���EÌ[t��I�Î @�3j!+�+ /әjҗ�2�ڻ�	�	`�-|�|ܲю���-%R�'F?OE4��Y��Q�*m��e�S�|J�LKa  C�]�ʆOUj>,Q&�!�s֕-[ޯ�]�Ys���5$]�^����7�y\ɪ0;����8m
	��L�e�t.3�7��LR)� �|4���З�z-�K���� �+r�'��]JaW��Rdb�8����1S%x�'8Z�Q���F�	}������R��ea��5�*𢅁&�Yw�.#�gE��H���{@��[%٭r�-R$�{�ե���t� �i��%��&�B�o�}6A�r�?P��s�Pϒ�8"�ލ�� ��u߷�՘�nn�"����!ޙf�KC_ZD�]<��`8�GC���ԩ��\���P��z��pBhm��Fi���X�붱Y8m������+��4�2��ق��z�����垇���5Q��wUFCA"�her��1rx�����$�$OHҊ}��.�X�6/wi�g�Y�]$�hU�.'�|+�;�����,ߛ��[��ZY���(g2\�X*#h��_��]��_��Q�/��Nl���\0���u2ݎ8S��`���w"=~�Vw�����_;	5��Pi4�U��f�8njY���i����@�Pg�L4�C� �dS�Kթ�Ѕ��逶da&���鮨�Et�y�w`����S� �Af���?H8���Rꊙ{^���4�^'E�f�p�HZ��v�[�Q�	f{=����KumȞҟ_�Q���.�&�;<Rl�;�.2�Krf�� �TLk�玻 )M����׻<˂^�'ϓn�ϐN�RO!fԲ�y�Z�����$���D�l43-� [�_�\,t�u�;K\Y��}�I���ՁC�a�S���#���%Uhg��<��yJ�f��ZpP��R1	�x=���w7�eVY���7��qn'o��4�$�:�PmE)�j�7Ԏ�4�mv}���>������zO$&�Ĩ]e��2��\�V��ɀ�D]��_B+��Q�[��9���ݑn���!]����3_�KZ��������^�S��(?�/�jHJI�P�2��������	��]����aa�w����`ζ�	䩛hY�.Y��1��k6@غ�O������z�J���k���'(��o�'T�	ص+��dw�SC\jLӋ��\;�0�>����y��������(��K'��@��(�Lg�*�g����
��us˃�MN��l�rR|�G�?M�5Fi^���b����ޢ@�����Խ���.�{��QK���ۋ"��ê��TB�h6`+ڇ[q���=)v�hJ��s�U+�#�q�P���5,Kq0�a�D�P���|����R
Hj�>���U�t���p2tEc��)dJ�+w�#�c�>�\�����L�F�t�W�����}$4���!	��"[�*}zs�=PH1b�B�.7���䥹��g�-n���첷�r[%v�059M���6��Sl��]��&�o�HF��Ҟ��q٦���V>($IF�:�B,1��+z浆M��������v�{�sPj�X�/�,�:D]��Dֳ��6^Ҷ�"m����<AƸ��j��k�3f1���7c�s��xG���t��G^PtY�n�+z�*�ó6��A\�i��/~��7T���^I�%.�弯
�c5���ݗx��2H��˶�ݮ�mZ��."UqwӬ�v�\�x ��6b/�Rxh��4���O���<�ȧ9�O]����X�&t$aQ�I>�\V5���_*�d9UV`����.�r��=Z�n��:i12��& ����Ⱦ��<tv�QM���W�W Bum��{��d�؟�D��5�p޶ô�E/[
Zfت6�9�&�֧vhT��W�v�bl�K1�b{Z�[oa����O��w?$�r�z������v��),#� ��0U�7Y�Q�(qs�ώ�-؆MCA'(.n5D
i��<��kǓQdo��ik�7�c W���� 1CZ�ݠ�f��3~�6�2����d�?��ʶ�*�I2����뿉T��/�M~�+�� a��z�g������@����v ���?�@��]��NEݾ�ƴe���G4$5N���c�D)�	
܁��~Ҽ2�&w\$~��Sx�Xh��5s;p?���_$��sk�̭kR<Os�{�c�^l3�bm��r�3�PXз�O��٬��mm�Z%%!���!�ObqN.�Բ�m�k,���94���I���PI�"���u�jw����U�I#�:J���@ՎP� ������7�W�tͮ���rC�߇�}9	��^r�����+�6����g�3w��%��3K�m+�'��D��'�0h��	�A���(^ڄ��;S�<�Jpy�\&7.8��Gx��b�$U�?Z�a?���,턪躢ΦA)xC�/�ۜ�I2CE5Й�M&�k����ٚ�x�� ,�&m�Cc̬�P#��Za�9\I���ϊz-������ ��x�
�^['W�a� ���WF����a��z�Fv�Q�ȦXQqΏ����qİ���홁h�"i{YQ��]Ay�8�>���3VP�
5R���M~}��l����ԅx`Y�H��"�Fi�W�L}H7s�,u%�+3%��(��XpЉ�i���Z�Ad9��RHx0N��p'�U�M7iJl���2MW^Aណ�G������tM-(��2������On���U,9�	r�2��5�y]���&�Sa;���7���C��?vk�H���A[=����*y�?�ʾ��j�(Dg��4�Q�a���-#�X�
��v�z��Mv(E������_P�Ûj>�x�{��P�{���u3�<ى�m��/H�!Bk����6�>��wP�[�P�К�J�����)hw�,�>A�g���C����ʯ٬eyddU~��U�|���#�ͭ"]�(���m�2�_^�R�W�A5���i ����8
��?��� &j�����r�T��Q�so�i���S4�nRP�@w���ˌ1}�����f���w�Xu�W��x��%����f�lxV�H��j֧	�T�up��3؝��G�0-�|b���\�����\F�or\Vh����,϶��C�xF/�}f�E[�3��:���I�`dX�@<"�,YȖ˥���dP�ԉ��SP���+��ޚG�����������G��GN�����Z,w�i��Oew��|Y�Ad��n�åI���1!"m)�9PG�A]�u"dL&�J�Hev��Ѣ���u���u=M���K��,M��h3}2: �ʣiu?u���W&2��X
�#d��'W�Cɩ��4��?���
#9������,��<�.��Ѣ�3���Ow� gCK�r��֏ޗ�s� �x�4�S��
�B(�M���﫪�qg�*݈-QR�[��,�?ʏ>vg�:�}YOn���,�g�S�ί%Y�$=4%�P?�4DY.b`�C���溘�`<7�Z�Yj+�eL���e��1˒h���D0�� ȞE���`fT�}=9�o$x�D����E	�6�?Rֵ��c���=������L^����]m���7H���
C��ś�8g�=���/Q�b<L��#=J( v娛@*>����4�Kp�q=���H�z�/�*�u6�(�\��d%oD@��(#�9W��Q++��L����c�����_c�`d�a�����ڴ#���G�kM���_��&f
m�-	�;9��)3֮JM᳴=b�l�����#[�0Ř00ͧ2�+��QK�Θ-�Uj�#Pݛ���6~�%�\�:�0ܜ��̼�]�^ /v�akb�!
����D�AK����O);�|R�g ����@ -�Ͷ
QD��R*�H�2|*!yUe�G)�z\$'���Ru���B�Ҏ�m=\���@)&�pDfD��'���Y������Z\���3�9Du���G�v�{j�`p� 1��>�f��p�b{�R�x���&��Ƞۙ��%AX��0��@�'AU�u�� ���Fc��P��>l�k,DQّ�|����O���Xc�/��W҈^�rdh�����Fߜ�x��I�����0kk�s��
��P�Xֺax�$��D����C��"���mW��	0H�����x>���,AL%�o,H4��B������X�-iǨd�IT.�x�p�OuW${ڼ�G����@��C1�@EO�F�n�`��e4NZΡ�Q߾~P�H(��	�NH]Z'x��O�����rh_1�f����$:�M����<ŕ��������f��Ъ�	L�rwE��þ-��}���)�o�Cx�+=l5�Mm+ �+���{�:?�XO�	g&���K|��~븊o�;��m����o#�	��_����F�h���~6hݎ�B�+��^��l���6�r���eƂ^�hm{`���M�qqIQ����#������94z.^�Cx�E¹��#��y�� r!=Bavwn_Κ_�8Y�9V����-�x�Q6�z �1.~b�HA��4ܭ"���@;���N?���� lC�nWQчΠ�>|o��Ms䲻ds�\��^���I���U�ʻ=�d�ff���/���\h�\CW(.n�G2�h����'�q�l���"�s6B\-u}�� y�1��fF��q1��k_�c$�L��i,�1�)����ܱ��N*�o��'�i'/�+�>ٮ58�����s�K���9�TS�jݒ��%�V�,�~�h�yQ~�c�4��Y�g���8��w �O}"<Y#�λ0S�ƇO2ɍ� ������X�$g���UpY��*{�ckv���@É'e��= �t?[�!�l�S�q|�ޚ'�~7�K��Pɂt�$Lx$D:s�>��}L�0�I����i�D췬��KHF��de��OĿ�~�,ލ0��l�-<3&�҉���iQ]�h#�Gz�e|q��J$��e��~�JV��8gDA�V|���{�+Z���/VƮ(���;{hֺ�BC��uTg����@�;�!`Ph�q4�N[�²�8p2-��3e%���w��t|���{T�d��	�I@fT�s�H	�ё���wބ�[�@dd*e�H?sn����P_��;��D���a�UM���)7M�
R�yW�t��X�P���� 1�E���5)�&9B�J�
�@�1�υ�K�NWfB�a����y�o}f4i�-��W�$GBDPC�E6V��Sr�_k�~�E&���?��pk%����v�;pN�R�E����?��~�?��5�a'<���ׁ�i�N|�!f�@ԨӼT�m�2C5����鐌t�EǞ�:>\�U�|[pЮ�> ��8ۏo,q8i�I%Gd�M�,���T���}p��c�rqp�h�A�	�_ �>���X�]��׋a�*�`n�I�Iv왡���7���G��`(*��IA3�&O�ZST��=P�dJu �鞻B��K��gy�m�Z����v�s�?iw�\�({�r��=|�Y�7���	/�
�v�\s��
��T������A�ܩ8-�B$���0|q�y�L1�m�g5]y"
�NG�gs�n�O�Q5�eJ�f��3.�w��.W�nc2 �z�:�=��m���p���]t�idhѰ :ٍ�Y��h��=!��3��͊/����SOa�z���>�[�3�o��N�0��S��M�X�߳����V�^��8�Q�[��Zٕ�5� I5���nOקS���d�E�����c+sZa�������]7�t�N?�W�6����Xc?A/_ֲj���^F1 ��Qٔ�M����[�}������N���[,O6WW��g��S
r��_f-��ڴ����$��B?�)�e Q�;%�S�^�x����#1fE�0Bo���z5���������H:Cj��򑕉��f��Oָz�����%~M�k�&��#����;�x3)ʭ��m�))��&6�|{��]��?ɷ�#\�u���(��`d.����4��.��@�!f~o����im�c���啻��б��j� ������d��5�R�u�z���u� ��yԍ$�h��;�1�ư���ώ��1uk}�͎%{�ܑ�/��Yw>�K�Wq���
�ւ7Ot�5��x-����:���(&�Fɋ��g_h8CLq�?9���|P�!t����B*ʕQ������>G��f˓�TE�6�&_v��b�W�9�t�����>�i�B����nM������{F���HD�t;�e'��p���Rf|枫h����qS@m�u���?qܢ��(0�u��l0b�D�ۨ�I���So�~�� 5����hok-J4%�r�վz��rz��=�'���,�p?�� LaI���If	=��S�x�]�Q��Yp�IH(�5�=D.Ŧ8y���Ydo��v�_���2���72t����J(�@Iv}{�Ѥz�^��iL����Q�QRJ�|����ȌP����_���3i���2�	%�}W��e��n��K���@h+��P���}��8S9�+�e-�=�l��ΚSd,�/�����b`���q�+-S�Q�ŬI�u`O���h�4�^��.�;��Ր���*���nMQE��5��IW$�N+�Zu4]�|rL�ܵ�b�����!��,�z�pew�lm�&���U����Q'��'2�rxㄪ2Ni�Aq5S����VdR�V���!��+T�~@3�2���6"��pJ�E"�3�����Y�M����QNM�T·T�l�G0�:�%Jb̚�� �l�,�>q��g�쮱��dW]���,��S\F�g����<�l�d��/㽽i+�Yݟ_�8�o���%f@�}7��"�xI;#�\�B�mf���o��g�D�Y��H���)N�ӟٟ��
־����%ޭ�晛OYt9F4���)AV3����0n���q���f��=��&�C2������W1�	�!��J��"��pK#h��aI�^�G88���ЮlG��J���L����}���#j��iK܋�3����J^�b}ļ3}�����/��Ξ�E��E�cc�����/!�VU)xzc'��I�|U�	���
p˳2sX��+5�uv�p,/�⤘�~-�������\�����y�u��98ܹ�H��n�%4�U��){��}��^��V�jPL�`��l��+O�O{����x�e1j�+/���2��u8� 4��7�}��3�QR��Хg:��5	o1R$q��z���`�Rqح��q�.�(ͩ��0��Kg%F��b��O���v�0�1<�Ruv�ؠ��AHY�hw3� h�$��g��U`?���=��q���Pl�V�~�9�BjK���P�&6�Ԁ�6Ei�5����鷳s�yHN���� [�g��фq�R���UyXlxV64EB     aca     2d0�9�Î�x�b�IjX��?��L�'�l� z�LX�a/�4���zh�%i`���_��4��zE.��li����OԲr�v_߁�W>\-{܊�r�,Ů�(Z�/7b�7�7W�_O�F���F=��9�J���W�2��9�!Q��	Ef��d��jDe``���Yͩɞ�ܶP$��I��V�U�i^6��v�C�e]������H�>6�����˯�>�v.lB�dh��h�2z�? 9�P�X�fо{`)S1�d��y�{)����<�UNЏ6]��*�tޫ���D�"8���� ���qh��⨆I��R��Dƺ*Vr�R72vL�f��͆r��$��X=��a%T�L�Y��[���ٖ�h�� yp�t��D�'��o�N��4�Z��a} �=���p��5�x��Q?���ܲ�&���[k��̡?����K�1Sr��]=�.̈�ݛ����O@�6G�h�K� eV\���3A��OP�m#��g���e�o�&Q=�~��19wZ��v���'���j���������4�6-&��;2��@��5U黁�[�o&��.V��z�0�,�C��Sđx��$h�y��,5����'��V�����7�s)�Ɣ������>�Ӽ��ǣ�c���"�~�9V%P���N��\��n0�r�[󟈐(�aH�Z��J����0#�H��
xE:G�;v�W�����I�7