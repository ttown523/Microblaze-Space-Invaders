XlxV64EB    15c4     850"b��ҁXc�D�x�۽A$l�e}I��Y���ȕT�� ��HDY��Ni'���(��6O��|�||D�����K��j�P/�M����>Iس]'�++�<���ad�/���1ڍhll6��515眧���y:�w��U*��=�GU��"�kmaΤXEْb~���;X�̉?��r�n_�\@`}�|�wb7��:W�=�]
��X֡��?�a�Gs�%o������*{ Q�$�Ͱ�F$b�ґP��bN�K.;c�2��fG���/PN�C�����Q��}��6�_;!�����ev��
CS��O�pF�SΓ�c�W��ۨ�{�y	.���N�ຐ��xI�D��P3��q,6x�a	C�Z��"ts�6++ѽvˉ��-.f�L��,��U�ϻ�KQ�'Q�N�����f�̓,�i$�4�卼��Э����"ǩۮ:�F̿}��[� ��ؠ����BR5H�x��kI�oǦ��3	�$���c0��Z.'Z5X���0�FU�s�����Y�F9��ő�'�g.�u���g��6��U�����Bl�,4�]l]��
g��!�C�6a#z-���2{$#��7%��U��k�N4Nu�y�83!�����v�gbyGC���3�G6�8O�R�"T�i%��}J���0����U��eY)�dm���k��� U܅yו��*��g���&�����w��?��� SE�ERR�b��('[���l�2\!"O5��������Kbu�"8�%�̇�B�Jd����JzkB�K�x��_��=1���#2�e�����e�]����&֭�C����!�%�b�7R�5��\F�?�KٿC��Q��ȧiXXI�l�. ]@�?�Q��Y�~�hE�O�uN`�;c�e��~r�]��|�FV`:@�5�_�xvD��4�PD��JS6���%U.&k  ��	<(ڠо��q�&>c�+�`N�P�A5��b�^���	_'�y�ro�<�7��?x-�1��8&x�)TO�� ���&���Fd�l�|~?����C�v�t�Or�@t7�@�k�4���x��z_�D�"��ԫ$��ԡ$ⷝ3/O/F���td��K���1��O%��G?��.�t}�L��T��
8%���D�Q�k`!�1x�8����b7�	�%�������w�m l�	�r�5��n��Wl��-���	B9���P��
�!�؀ԍ���P��m��®���	�j�e5x$zWmB[��OP,in�Wt��Rޠ���J|M�ұ�3o�c�hzc���X����L�IRgm�틒�o����g�:�9J�b.�0p����R�1��d������̠Nv����p��$�����k b�ԗ\ٕտt��ͳzǋ�+ۗT3ҫ���5N()Q�#�~�Z~ϧ�2ogN��}i%�n��*����ej�xm-͠C���ekG�?����>���o�8&�;8��v��m$2��&��������ܺ�bQ���f�څ�mIE��S�}�˼V/�rvv�Ȍ����Xn���߸B+����ձ g�Mu��q�M����օN��"��:-R �����#?���'��3<ڏ���j4�T�M�z�������إ�ĶJ?�����Tɂ�ľ[|@:��R����d?���%��.�҇�45�,f��/�0Z�i���߻ۻ���{�hE��bǳZ�ˠ�x^9��1wb�֠
�c9��ru����l�a_��Pq���X{���J/�滉[	m���o�,L�Yت���H�#����z�u�RI����qV"gX_�k����W¬,hQ��Ӥ	�V3ҙ%�!�Z���u�#դ�2K^��m�o$�3����v�����eV��Z]6�C����G�ꊪj�D���t�D�H��3i�!3�űf0K���WXbG�<��LO��#pd��~YH�q���4V��m�du�;IL=�.�
xc5M�W��t����U�8�3���į�3��TN�.�eRm�2�\#�뀘E
 �ze���ȡs�v�|�8����O�L���TT�������#9�˗~�/Ya�