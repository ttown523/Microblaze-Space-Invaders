XlxV64EB    fa00    2ee00H%�_��P:p���F�׵�I��~~��Z;��K]��ε��`x�Xo��{���3�%ai^�,N#4�o@��Gڣ�+��r��'�~�t���-����f��O��g�����mw�sH��OhzlX|�Z�6��x�EЩ������G���pe��l~߳��P��3r�O���e���J�I�u���J���U��o�e�U7���d%�Q�<�%t�{2�/�e�!�NXJ�g3�-^{����{r�;i�K%�c�S����coV�Q��a�xCi@� �y^�𼡔�6�),�:�p����J&P�`԰��ߗ���9�]Iר�U�V-�ds�S	�(�HѨ�wWg��0r7�6N�G[�W�N=�6��n�������4�;}EC]�DO���}��b��6h��AZ����'Uk�I�P<���!+�D���R¤7����Քj�ӊU��ɿ��4"���Q���r7�6�L���h�������[t?0�ʩ�N�Վ��~B6븖�a�50W���w)�^A����{��gH�H}����B��k���8Px�!�Bg�!��b�e�|���6�ն�h����=�z����LG	x�2x� X2c��E���a�M��F�Q���5���[kN��n�� �A�]~�H�t����r���#�@���[aG�uF%yvB��+ۄ ���tR[�T�̼(��o�%{��z�k�p���uT�� �L�}��C�L��@
k��=�d��BQ��+�E���� 4V[�F4����,�D8�)1̶7���mqF�n��{6Q��V*$��qׁf�1�,��T�%*�Q�f�ݯ����?�����l���#�D����(X������T��W��i.-�Z��傫� z��03n|N:p�	�Z}@#b��RM���Z���f��
	?��`)e�����:���:�%�����䭟��<�D��-i�x}�*�g[qZQm@��d� �J���b�u�������W�9*k���A���f?���&r��`��C�/��"�j�n�^=%��+o�ß��R���	�6�"4���=���lR��o�n�FĠD酕I�v6�鋪���5Y��\p� �h
#n(�G��jqC�o��E��D)~G�4	g�V^;�w0�D}�S�o6>����.0��IH��+��t[4&ˡ��':��ڐ��P�ӟ���PV`*�ԯ<��ՙ㟼a�U��X���s�pV%��,l�Ib��)?��]^%���j<�oPF�GD�!:Ehڥau i�cl�������!��`����\^�k��(Gp��t���
�1�{k���l.�)��ߛ�]�hT�����m�!��1�]-vs��v�!�_J�ä�ѧ�i�L�����LQǕ�Q�a"��k��ݔ*TUK��J)�p�������Q�PD�e�6c��r��z����K�!�.7�;xv#���X
��G�τf�Qf぀���]�g������<�<�+���<�h��yp,}�N�z9��@V��^� P�@��h���d5饷��g��x��0�k)�[�3�8�i����� 3�@:)|#���a^��rM�ѵ�����h��%�hV|a�t��ǎ2;����ت9x�J�}Z�HSV�j���M���8���Ȣ��!�'����=����:�uƩh��^��)E�t�i��v�����WV|*v�s1�[�'=����}C3`��;κҢ3�����n�y�Vxl��
�OL�����uQG �_��ؔMg��a�C��wè̔�5�ÏQN-r��ή�ݨ\R�OM�%�lVaq��tx���4��N�ys����?�V��X�O���"g�候Z�q(6R�-��Ȉ���u���"��]���te��3����� ��/��1DEO��{2d� �Hx�ZՉ	I�{�֔��S�~�^-$�!�x�R��J (�?��2�v�'E?���t���J�0;da�����T��w���/'� ��|���\6��ol��e�7��I��q���k������~y�P<x6��p8�͙A�t���^����C<�^�F�S/V��*F�'�;sa��.g��Ȟb��U�����g��&HV�/����lk~�$����$/N�&���>��߉�&7��%�{�x���˰w�����jc˱�����y�Y��IJ'h���}&�����sWd)a�b�s�AN�2�	?�_��
|DD��(�,���8=�묠S-4 %�?�����j9��g�HU����߿�Q��D?L��(�iTsr2�a��oL�"Mv�$��6L]���^��%l���i���=O=.��֨��GN�Eٞ[�����I�vޠ`�G������*"+h��w�A:=q�0�g�}��R{D���{��f�&���9|�nӢN���z^���#\�J^}z&�8[�|V�R�c��ӵ���6e����\O���X%[��.��=��0*��')����־���Z1h����J}�<r�' !��E���Iqf�7x`����� ̼r��[�W	?���/(Ъįd>'ŵf��cԫ��d�d�	�rL�a�Wf��At57e�,��M�&�~q��{v�T�i����XG�8���j>�{ݥ�pS2�T1�=˅�
$�L*�f\���g�J�=H��>�tx��S���� ��E��?q`�J#j��͵w@�X%"	�s����)=J-�����
1<�I�����Lr�!U5��$���iX��d��R�_s*���ߺM��tz�<�	I���?�fG!p=h������4r,���6J]k"$v�\�=�w(�B��¯�n<����I�]#��-	}�������ho��ބx�f�(��ځ�}�g��n�>���}�(vr�"�:�L�&����*��-���=�o9�R�~�0�P�Y�)A�|{�����v�yTwm)<V9k.�
Vla|�O%��rh`�7G�mW�����W��
8F�,�H��W�X�\&��"y�ժ�Ƣ'%>T��Nj\l�q��}�j0�k��!���qV���F���A�D�+����SL8�D�����Ȓ?W�8H�]`�qU�E�Ǫݠ'ڠ��^�v6LA�)����EuUn�c�W��E�Oi�T=u�x��z�Џ����Æ�PW
�餪��-*�(?���9t~��&
�Z�IW� �m�ǥ�α�\,��9��IG4ҚhX H��t^�l�٦R���J�������n)��r���,���T�q쓐�S���U`X��F��]T��㮬�6TQ�	p����&�h��@�IF�œ1����hP�f�A)<K��M{�t�$�A�1M�T�r���^�,3�v!x�8�5��ya�
����'��M���Te�@��[�[��+�~����'36�m��-q r�Rk6�6��?7P�4�1cɭ�-�����������	+Oj�g�UU�Ҥ&(�_����y1���RM��;ݼ���Qv����˗9����A*t,��Q�H��IO�7b�j��c h˲�O�q�{����i59�6d�-d��B1j�����>�Q�5�Pq����#M�|C:�\�����R���
�7�?}�^�;{R-.n��yA�D�Ʒ*���h�/&��/��y"�v�r�ۖO�w��3TR���_��C-�+��"Ƚ2>���;��ڭI�>s�WWc�n�D�j�h��T�GQV�d�N�#�7m��;�΋iK�����sc���Y�J�����z�5g�W|tǐ��;ݢLz^oq�	'|��� w%Zsx�Do�#��!L��*�%u�ǨN�F
uŢ&h"���"���c�������;?� ]K5PnkH���S<��hvE�+~�בe����h��#G�C��b���&��&�R.�d�w`7��m[��`!��8���R7�1e�>��ɫ>@'F�(z�C�}�.@!>�8O�2���F���	$�R��z��t:�>�Z�_$&���22�,��̋ZR��B*����:5-څ���,��B�;���z�|D&&8;B�{'��˴�C56=9z����V#:/f���C)9�B&c��h����Z�Ӧ��$0���q���m���7�$�mы,{��5+�T/0�u�7��	s4�a�Q��Eb��7�b�f��: w�E�dֵYm,lJhR��]���F�zצ'&r1�"=�:O��<~e?�|��s�7�פ����ŋ�џ @��r_{��թ�K͖�fGvC��,��2�M1,�o��M�?*��*x���{�8�of�4g���E�@�o����r�[�@ռ.�^�ܯ�c�xץ���� ��&��O��@���v�%n� ���7؅P�n��j�`{�E!�$���/����)X⑂���i�@<"��J���Ƀ�\B�؜���[��Z���u|���'_U��|��@���W�O6`7�kD4����/�+��ZC�N��8�	.���?�^B����v��n��E�ƂW�̲fF-AB� ~k`�c�C�s���z�g���.`
2�$�E��)�\���8%����x4<ƪ��i�(��4� k��Hwk!q��um�X6D��J��3�&�UA�[?�*֬�͇!H@n�ؐ�y3~C��͠XB����uoO㟿����VIh��0g�x��`�+դ�H<O˱X�=OB��/���������B�����86=ʉ���ʤ��:ցYJa�j���h�yrF=�@��x���R`�bh����0���ڼ�����5��~5���ۆ�`'�zY@bTJ��́km��]�4���o>4�����Qe�����bU;�.~LK��.��=H��.&�T@&�ag�-�i�ޜ#�H�@�� e�'�":YT*����2��آ�>���;�T��<������c|���V~ް��0���f�0\����|��Fg
tعI"?T�D����d�%�L���]��T0(+!����xHeU�]OOI?q��i"E��f�B�MQ �N����J�|��ceR{�=�7���z�� ��b����Q⳹y��l���~�̬ٹ��YCZ&��hg+?�k�Y��v�t�ˏzj�d��_6����_�]kj]]�7�����;u���;9>�F`����BT����	��<٩4gLyk�Z��jROS�Kl1��4*=�E�iY�;�~o�[g	��Ci\?�o��e�ܼ�1�i\����#Q�U0 ��X�$Sk�������[>�"ԼWc����_a�����ߣUb�Hb�q&@­��j?��99$��!Q��b�R�������r�)�-4�jЊZD��I� �~����sa�9�����s�.Oq�i+3�wqY��6�Rh���T�*���zu�Bdc�ޓ,�(�Q"[uj{���'�SY.!�6 Α��~�ߚ9�(�֭4�"ő�bO�l85��#�(���E�����;��xBY3�p�����~��
��B��]��#��8p޹=�aZ8��0eX�e?4蔕����qe��в��s0���#ȂҞ��%|���:���@���P���8��`4�A��n"k�`Ts2o�ɺ_ \$�iݐ���ZdRjE�l����}(0��XM%s�������\��!�[�ϛ�⹋v;&fk]�p�{��_���M	��+�Zc\R�E�]�TZ�$4s��QWs�/���I���L��U�e�� ^�-�a�|�i^��QTd���R���m)鮦n�{/
)�ȇ��O�5���ﰭ�3)�F�o�|��@�%$�fsZ�	H�t�?}���.w��rf۠/�Ϯ��gn>����&�Νv�ߧ�²�d�w��D}pm�v��� �d'��aU1-͇O��f?�W8��Fɝ	z��=������)�c
L���l�������$x��� ,7Ǎ6���d��o�]*��)�φ�4�oV�Ny� �����,�c�G��p���L�{{���.M�į�h� Ź��t�`wGo��9�j�@�~�
)���(����7���[O\�>ZI��702�؅��Y���q�Z};���$���������������SZ��P֗p��#���Z(R-g��@?��h«�%c���q�Q��v/&��o���ߒ���(\��-����ۛ���U,zwօ&�?_v��r���8�M�,-�9/XRDwʻh��:~�$���4j���+�����}�n�~n����خx���;�^�����f�>7��%q��d���~`��B0��1���}�M{^���HIv����(k1"��@Ĕ ϭ�����)�}���}�#;`"�!�f|���/x�b��9U�4�@�����<�2d����t`T_=l�\��-����)އ8x$�{'�,���:�ځ1�Z�;j��Z���:��ׁ_;b}S�m`��1�oyU�4��"`�6�$_���J����W5����tYJځ[���n͹��{�-��|g��}�3?���a�囒HN�O��W�smw�����W�=zt�_]n=�+��֎F�6/ӎ؇���a�| �hԲ��Fٮ���]����ʘ�#���=�8*�5��Gdq��e�L?�J�:/,k�gcX�����&n���:��OkiES�O)���֝�87���9�9	R�3�S/�!T�.��e���C;�;�V�k�䀪Q�g�Op6��V���˩V!KϖM�jt Zy'�!��h�d,rA��%l��|F��8�˟p��Xb�]������ѐ�o􎊜̣U̲�u{?�<���(��n�	��n�8,�#��<`���vhR������d%��� l��PZ�ϽJ3
����8o�'1�dw�](�:�M�\v����
 ���A�>��n%5��C�[_
VЇ�v�g/��?m��k��E���@v��ID^h[\��x��q�+����ȲBƐ��(���F�.��d%��v;�$��A�ڥ}�@ً�u�zs��0�*�D�Dլ�s��Қ�m%9���Ώ�N�+��v}�b�lnƔn�J�;	w�M��H�򿰘����]�^)ک���I5�n1�Sw�������P�ʚn�b�.t��=��m���SV���?��ϫ�l_�ܸ�=XϕV
u���L2A  *���q�x�p��
�ךY��N�
l���ߛ�U��DZ}��ea�?7��/uMXO��BV1ް����:ܻ�+}��k��8�(.�s �;4h_�rېx$_��������*nP;A=�<u����(�<�q a���H֮yc�9���	��w4��P�YH�[��ngj1�g�ڕ��r�nX+�G���������Ԁ�}��R��
6���T!2���PE�4�ӝ�`Iڟ��Cq�"��K`7 lNj:7p�o{��޶�_���LȠ��d0B�oj�R�F$�2An�q�d��a%BءY�,M�����3N�D@o�h��%y:Fg�2�1,-�Syg�Vm��b���b9�`�D$�^@��]��mS���٭�lLO���t�K�¯DN���C��#m�p��xy����K�dv�M:��R��	H@���r�#F������Y����G	+B������X�F�X��Œ���w�0;�^<`��\�!��x�Q�*�r8'���9v�:���$���yo�=�A��,�Ur���
�#���IH�Z�r� <u"�[ɭb9���1��$a�����㊩|�v��δ�tr�m�X(o\������Sl^�xwٶߋ�8,�`���Qu�����&��o��hnrZ��q>� �i 5�'���%���=Mø��:q�p	�:�p;��D��4����
�#E���@|:���h�"3�Zsm� )��#�۩y<��6?�����a��cOt"��d���/�CS=���R����H��Ir��[ Tnc��B4 ��ZWf����/�w�y���g�:�`1sٴ���$����̺�Rh�������"�]�4��K��A�Q|b�6)VcK~�q)A���<t��Ē��u�ˑ���"<G�\��� J�ޘ���˪x�vQ�D�nh���8{��܉��%
�
����4�n�~�:خ�����*�IC�M�MY������:β���w��Y#�jGDŰGa��f�|(�s�`������f�Q>.��/���D�:�B��x�gS8�{�O�[�Y��2Ůo�D���JD)�f�$BH{��{�b���"4I�T;��ћ�H����� &C��Wh��O�:iE�̬��m㧶\���8>Q�{�kC9��2=<a?�'�;�! ��Eb��үDp� �r����2(k-�
�Ӕ���ɯ�F���e �v]�_|�͝)F]l;�8eH�@���2*<�^��"W��-)�������L�}�f�\;/Et���,s���%����p�-=6��6P�S��e5���ey�|��v,G�uza��(Hb�b�Y���E�,���-�u~u�j9�4�ц\���CfCn[�&i���^kL���T`�����$����?��2�N	�#�b!=�ah�m|�4�XAu%Ze�Z����9�v�v��{1���Pqu\e櫉\�ciFW:u@V�C�
�~6QC����ї�z��ly<_1��P���ա�q߽�u��d>v1u�TӇ��ԍur�����[�|�خ���?N������:ȘC&��4��9:s��Ҿ@��՛��J��+m\�ྲྀ�=|P�Ki�a�ǆD���z���f_ࡢb���jRmY ��2��IqI�� �Gfct�����7��S/�08�S!�y:ܞq"��LĴ���*��=����*�d��A������S�����Vhh��H�`R�
��Ľ=:y��@b�3�Q�_ߪ�{�{	=��r^��ɪ�KU��ʆⴟs�s|-����9P�(�z-,��� ���m�@Y�M,4�A��Il!r",:}�yqF+��{����*�6{�[���rr;��c��8�G�A�����ۇ ���<5o�1�h�2�
jR��]���p��Q�rE0��3ƭ�`���_��5R'*g�ݜ��a m����w"�-'[��4�Z�H�=*i�}dЍI'����k1z�6��3+�9$yQl� ��_!7���@�>��4]J�M�1B(�����:�x�	U��+ơ����={Y{�d9�������r�tn����٠~[ŕ��_��aHD4�bV(Fxv�@^�&�N���zL|��O^}��$�f[^���DIo�n>��D�M�}�F�1s�Ц�pff�Q�Z�o��,�7�����!��Q�n/K���G�Lf8� Q�M*߰�����X-��_3_jK�<�Mݔ:r�N1H��8Uz��áf(<n��ck��M���SYR/i�Y-Ŝ�{$8�*Ѳv��2�w|&���)e��޴���^���"�Ч�/S"����n�CPÚ�\$4ZXeTXQm}�|�F1`�`<s����N��<�RZDqTw�Ѥ��
�qOC{|��(�W��C��~�$�z�!	D�����G���� �� �٢�M�\��f��e��xo��ç�(=�N���h�Ψ�GP���)��o��>ȴT����gM�������&� �Yl2q��N%�*W��]�+�1�j��N�<��i�t�r#�>��Pd�݌_~�����X�*^DEP:��ߡ�d��w?�$"}�wX��� ����G;O:��<���4}�f.e�ښ{ �޼o6�	-B�48���K�)���o�ˬ�s!���9����o��U!�����'�4�ǽ�K��U w�/�
���~Z��L�JdlbmvB��I���4ɲs��>6Ϫxn��9O�w�?׻V��]�?�r挿m�#c�W,�Q�k�?�gM���'���9?[�n����~6>��Eɪ� k���.�,��>�W�2P�j���;�*%�@�vz$��#YWGEU����ȧ�Id�B�q˩[���d�����{�5�_� A����-�t�j��q�28�әm�77���W���	:7����x�.�Cl�]?��M�Ni��{JUS&W-�����u:9��@t��$ Џ�7�<��CEUh�<҂�C�Dx�=�`��{��'~��b?�ӷ� �q�(�7�n�l�۔۱�TLEb���V����	Ӿi򼟼���%�� ;V�_F�w�>u�n���� a�y*E��lM�i/�����x�5ׁ�i��h/cO����2�bç_��Q���7٪��Hz`aX`w X�;�{+ ��D���T8x�Ƨ@�ۧ6�NP���r�����<�ėI��	�"�U�h����4�����9q�Eڀ���Ӗ��Lk痳�,�%BcФE+S���]k^���y��8�S�ܵՐ�� +�*������gT��~e�c�zU��� <
�ϻ�Z�IE���)\6��k�p���G6�����ɛ��iUz�R؏�?���<߯�,�&��v��)��5�x��ҏ�;AA~3��a�a��	�ͨ򜾥�Z,~T�*���>��خ@yg��o���6��8���uJh�#j�5���H��\۾M��'v�e@�9Z� �kQD��P�nO��i�u�}�&.���M!y��D����0I�0#�!�a���+ǵ�g�8�0��S��~(�����/喪Q�}�����(�*������:6O����G�=�S�(¦��C"e�L��>��JŜM��j|���V�]�R��s��NF���'̴������p�S1z;(���B�X�v�T�[�9�+��<��N���O�k�J��~�ٞ�a3��j	���=���hA���42��x�R-»�ow�t��7�K��aSv�"~�0Rb��鉈@ _�8nYUE��CP�;)Ȧw#e�L��M��k��Ňa�TLY�ke�`E�����U*�	�A9L��4Z��/�I�ZY�2�F5#l��<�w--�qqφW���1�/�*ف�ʉ�q]���R)j�<�p��n��}z��Z��@�1��^o_1��X��#�%J����G�.��12@$��?=>�L�9��}i�6��@'][��VP���`#޾T4�c��"a��t���l���\�E��,!kBm�uv��B��A��[���Н,�k����_�1!*���%'��y����c�-g7R�#�����K#����J�-��[�{�ǯ��E��g1:����Y�:�M�Қ��g[q[V�sBs_F��BO��7��j���#�N `7Pl��|%�O-����}�$�(z���C�X����&���6��4=��4����Dt�9������<�}�n(=rq�����Z��ЭqL[�ȇǮ�ǙN&�����Ǒ��Ж��F����K�Ζw����u����P%�ZSf���w{䤵*ފ���?(0-a��V�)e;�b�-4��tf���$q͕�\�#v�t���D�N�R�'��RF�$�_9<�9�|��0���V<�Ñ�)�u҆�;:d/��A��m�$�y����=�rzT��)dI<Y��E�b�8�>vz�ʒ��
#5@�y+u�
��y}AVI'yx�%��q���m�?]��쎼0U����$W��>FFN�.���a���N����}l�s��F�C7��f���LUǉ�q'a��)�M�|��;F�V�qrbc�=.,D���ܹx��}�5ԝn~5#k؟t���BTQ��ۨ����5Z҇����.1kJ��M5�\��]�ʈ�Օg�E�Lj3�����^�].�}F��XlxV64EB    fa00    2c50~��3�n qԽ!j�o�'��^c�^ ��99�d0X%r�:��ęt;|b�"Z��2�a#f$��#\�h֒��P/���#BUj����*<�ە��D�OlS�~�"�tv<�W��h_F���k}S�HlhS�U�O�������u���3���LM�_��&z|�i������ϩ��H����+�D��]q�c���˒�#���4�	�okuύN'3�1��adS�@��~{�ڕ��nO5�˩Z]�r0��e�gTUu��)��3�����vB�e#J $���v[��-�G���o?�
s�Z�~�NST��L:��=�(b��4�l1�N{R���5��M������p>|E�Ii���Ѕ4G\N��ک}���Ⱥ�Fg�5��ڬ׳��/סV����2����C��z��O'�5����,���Zh�p{����S)K�F՚�>Y0#R��B��u�(F�/�ơ"{�h0��H�
:����MM?�qj�������q�)e�M�E��6�]���(d���4���� }��k�-V=�9��0�]�*���!�z3t��1Uy�i����ޔ}��4l!�>e�80H��n��G�3����[��Wb��9�p�26��km۲��2�������(���G���6�/�/j#�u�bU�z`�2b>�=�(�Ut�H�FO�{�:)}En������q�C� n�y��Z������|���9���^�q�7��������)���O\E#_�1�g�w7	��0�orL�"DF�68:�S�H��X��u�O��Pi�8U��O���q�p��x�+�n��
��u/�T�u�,!���|�5�%�c�x����X��e�lw;a�X��\�W�2b	y҃��#6b��E@;��	Q�=�����'��yi���B��t�Y��D$cw�T��A��]m���߅!�BT�j1�tx���e.6#�ﮛT�1�k:���Z?��}Xf)�R����ݏ-�B:�����w� Y-Td�1��ĺU�Tգ�����B��s�|"�.�Z���R��.w��B{�>}��^%Md��Čuψ�m�
�N�d��9��F�g�������j�W��n���O��$*�!�be�㋾Z#�<�ʮz+��fp�ll���1lt$>�rӘG3��ѩ�>rAE�FnT8�f���-�!هQW�9Rt�^�K�Nb=�7n�	���Z��@G&��efJ�GuT:)�#@�������Ѩ&�n{ܩ�x��=��ț��mXigbW�w��:@>(U�j;���fzv5��C��NfN��Y�6��d��茙�X ��@i���+�XW%j�%���I����`����x� ��;��F"/MJ���e�!�Nn�����-j�]IS�,�m��ƅAzE���5��P�1��z1h�d�T�g��0�"�\K�;ǰ��/�s/j-0y�k�8��8����]3�S��!3�1���n����=�X���~k14�f��6Gn>t{��]���s�7�y% ��P����0�k��9��"�"Pa�-��Z��k�>� �&��}���ц��쟉`	���C���Z}$�ฑ�F����c���o�ph�Kz�(%�]���`fz씟e���7�Ͷ̈́�����<� �RL�(��?-�A��LF�
����B�QG��PUg�7���A��cqwI���b�*G-0��.I�~�.���<�������������GmÆ��ʟٙfM��>����}t���yŐ���T�T�q���ipԟ�	�r��74�`��//I�`A(�d�a��Z���i*�ۢ1]������L�����p[)�y�p�G23���Gض�D�}��]��h�\9܄ř`z��6���fG�B\��w��_�ʓU%�� �Êq�]ODu���!�b��~4 �Q���4R� �p�(:x)�t�'�����P��A��:�"���p�P�^9�S�}d�@$�Lߏ.�d��mD�s���4��suѷ#5���x�_�V�Wx��r@M	�Ng�x��C��O�_M��)�{�ە�������s�z���yܥA:r�r�E�y~����iv�O�*a���a��V���MLG]�<�a������[Q~a0g�#��*h0�����.�&M�~ Ҽ\	�7��V���A���߶@��Ƿ����cǢ��*ƥ�M�;��ϣ��G���2���r+��J�kp2StE����Bw����[t�`T� ��P��fR��:-�)
//����][�r�K"�/������H�M�M�C��l�Z��,����� ��_�f΋�Ŋ����<��-���D�~Ba��T<�����ŀ�Ĕ+�Êi�6&n�2\NG�S�J"s���P��:c6��a�� ��_e��GP�bIZ���o&�+v
$(�/k`Bp����)j��Xǫ�hZ�3%�j�<���jN�e�!
�k\����!�k����#~g�"����=��U�̒�������VO(Hx�d�)?��5/�����yae ђ��
i���4�4�6s1,��QE��I�����T�h"Ns�2}�'��"����A�����r((C�H�/�+-ژ~�܈��y���)�u3ȟ��3C�Ė\���t�����6}K����_�i�\��%tX��+�5 ��au>��W� �ڭF�Ռ��d���,��s��<�����B�X�H�z�}Q�f�i%��Ip��Չ��`�%5X�
�g� �|`�*�����P^�X㸑��=z�P(�,����c��+,����ҫ��o�ұj<r_d����s,?o+`�!B�PL���!� �S#�VƋ����<!r߇n�У<���?e3���Ʈ���K�;H�\TM�J
�,�+���i�-N�k��爻��K��zj�6�[��I=�V�	���>Cݰm =�7j�A����_b���H]�+�|vْ�����BI�I�MJe����06�
�������� �T�YD��!�i�E�	Q���J�G2P9@]| Ux�2M�#�0�|��S'H}������r��0�DhJSa.p� ����H�����=��5!:oΌB���4h8Z��VR3=G\'�[��+�Aen�y��8m��wW���κj�8w~T;���QU5�x���v���b0[r��rC?�(i�D	n����`K?ٹ�q��G�(d]�����B��#�$zr�3�S�Y~o�]�0f���Ͳ����ٯ�0��~D�'����uS������d��W`<XA�np�a[6��TV���~�}(��hby�����(;Tm�|����o�8�!*��y�7#�,M��9@�����U���5l1�xV�V���]HK�t�4�wO7ua�����I��ϰ|�Tі��*(:�w#���y�q5<N�vl\��H�lT�P$��pb��J�i�@���5�hx����q�!�����<�!~���~�Η�A�	��:�n��
�F�^��)?�3
�]��>S��֭E:5b�U�)�R�tU���j�Ƶt �x�k�N Ϟr��dM�9z&�z�v��y��e����QK�$�P�35��PuC�6��:�_��}��y�0���!��(?��P@���wr8��ӥ�1(}=zaR�\�_���FQ����0 ֞�|��>8�ؐ���0���1l�P<�]�>j.Ƕ�gԬ��{Hu����6ȋ��7����4[����_��R�@�����k׍��~���xC����4C����?\����gêA��Zy��7_TMT�׼Mku���:u� ��tM�H�~J�f�D�K@3�5����Q׊�B
j�asX��˫�tB.7�N�L�l�����/���k�Xa�zӧ��zҥc��r����4~YsV��V��v����s;��d'�����%���G塄8� I~o���
,G�[G��tX�G{Z�Ʊ��4}�s�q;AEm�ä�����ml|X�������-���#ΟQКv����MS�/�i��¡����!�3�g��m�1W-4��OW��6W$���E�c����� �N5���)��7�6i����O��u��^,�1}��iȨ;�ؒy��7׻4�Ԍh̮�]�&OM N��h�|0�/�~>5@d�xѢ�a�l:����J�4�����"�ڌ�2)֦/���,��G������~6fm��� �+��3������z��_w�Y�E���R�v�kE����K������@��]��Q;�d�zBQ����wp��쯜��5�=#�|nC+{���^�H�?���˾� c�GE����TZ�������,զx�Wĕ	��p|�6 U��x;8��y>uv�(b�<��o��dA��AOD�"S����rǾE�>��8�B��8ҥ�v�@\�9ð��iqH���֯ܡ��T8k��h�)ܬ޳�@��`i[^�i'� U!ӌ�`��Xm�0ɡ����Q랰;Yd�v	�K�J��x?C�����1N�-z� LM"���! ����SǮ9��it�ԩ��k��v~R'�5uV��ʇ�"1��o����a�tWvrh4�Q	��nI�Ŏ�A2u�X��=c���O>�e��x���.c���>\��z�,Z��AZf�i�b�F�&׭�ZA��-�P5S�I0٪.�Y�7���b=�`�GN���`'��_��e;�ʙ��!�v���c���M�l{��3c���0�[J7�>�q��C� ��`��G]�iR��W{��e�t_8�.�e�D��Tc��)З1��R�F]O�M�)w���
��\�[<-���a�����Ď�s������V�H����݄!*�`�b�<��|ܮ�ޖ.��:��-yd�0�s�Ҁ���/��h�y����aә�ĶoQlԘ�k/��Ɓ�������)+[ �||�?�jƈ#U2��K:�I�N���\]�,cj�SF����@5���f`��"4�ߖB������s�A������3�f���'�B�/�uk�q �_ ��f����)�4t�wa�Eq�?�x͝��ih�4kcK�!.�*�6�T���Y���R������G��U�G?�R/%�_.m��x�"=��.���9=!µ��O�y���lF�͢p��a��Q��0rf)�,��c*��Z嬋v*��"��#���T8 ���f#�:�u	)�̨�!s,#1��(�a��c��W���Y�*�A�Y��A�����?>DK���y^�������аn�OTAy��V�J�N�Pq�gNn�-n&�� Q���� ��L(-�%.;M�� F4�
 �,:��k!�_q ��΅�5��X�����Aj<����n%�6lw�hB�x��t +�����PI}_8����Q�§$�Y� ^Φ��߯�F�T`���c�CB���aU��7�ءȷ~����˷%ܗ6qI:Yt��qY(��;U,oʕ@ҟ��<ԦƎo��/�����O���C�;m)urd�[L\��_��d� gP��!�K1�*��=��_`�e#"���Ƀۨw=>��=��|%��ȻP�.P�z����F4q���fr7�CƄ��埩73�+T�eW�>  �
]h�?اUg�Iy^��i�l�o���"�^�@���� ��mS^f'2�%��0�|�kl�� �R��,���G��ژ����,e� �����S���nwf$)?~��N�9W-'w�v��x%V)��솽we���D�cIb�	�'�YS��J���B�-W�Dǒ$�����xC2�/���DC�e��3F#ם�|o�[� a����F�^C�4�i;��F���"�ẑ�NyV6>F�I��w�pL�|I"�-�^++�WH�{���n	b�κ����0��ǖ�c�y��.�(���+#�O��9���&�v��	Ƈ����;H��|�� �Aێe�����He�pN��\;J�f!͞�E����uΫ��g���s�"�\9 ,�Z�����<�YK��b��Ђ�tɓ�t�U�h�,�lz��Q���������9x�͸!�3���"���ِMp��I� @���؝�[��s�[p��"�Ť��cU@:�ǦH8f��m��wvdX���٩����a�
̫��x���Zo(?�[���+��QI��?�?�_����8�xٙ$�P��'2�9�Mi%Z!"Lχd���q�Z�������h\vohF<����?�D�;�����
��n�r-:���j}��\��e�Ԗ�	A��x���O�䊇�-8vh���d�n	~������q:?2�i
8�j���"�ڿ���HSz6G��ٱ�Y����ۡ>��cA,?q�ϻ�frb"��u���%A�ev�i���舔����ä&l��4ج	B:�q2/J��e��w 8Qw6��-#��/}e����Ĥ��jX�t��u�mG]�X'���N>k$ G���dS����ϩ��Ԯ�>��ˋ��F	׮Z�m]���wj�@���}��/zE�V���wr� =�!���&�b�Oa�q����Ƞ�;Q��
���h�q&u��,��|�t��̥���\Fjf��<�/d�n5K�7�����%n�8�V4�z���S����ο�1����Dߓ�;c���6��J�)�H��3˦��2?����JFdU�rǜF�,T&��EJ����Wo(����K���8Bb�IT����_��/<U�mI�7��:������k3#;�R���ЃK�����(DnF�<_�q�J����.���C��A~�JM�SE��x���G�n�Ty�I������4<�J?�����[ ߵ��"V�A���dD8��x|.��=zpo���?椅���B�Us�x�&��,�d��C���[T��]�Z}Kų�y_�?��wDr��!跅�揕�*OXu�j�x�g�k"��u�o� ;eQ�yEˎs���	�����ե�B�_BZ]hi�)J���� ���᳭��,��d$���u,��)򸬈o5e�O�"�\��
�C�q���D����o��;U��&.��O�%��}Q~�B����iA��y,��f׆�������FD4iePћV��+��-=�;7��q�Z������@��U�����Wp��0��1��Ô��/���7ܥ�cj�?2���K �(���A��N	u�L� N�a�ש���'r�4�o�������Jş�l^�Hb��"1�X@m��E��P�u?��ۣE��D뿍����z������/G� ��V��tۆ"c��vc:SE���9:�V��`V=���[���Nڶ�l�?ZYZ �0����[�`����#/V@P&�(�����+1]hC.9���~%����3Wp���9����x�O�|�yu[ =ð��)U�Q��b��>�zy�i+YLN���an�Fs��:r��1������������;Z16c_�U>��$b1�^
�{=-�cȹtKx�^�|�Ǘo��U\����\�4��Vc�МbnjL�/n�Ӣ����s^����1/�9	c�A�X��Mfߎ�O ��#-�枆�}4�E	1E��~�P����o�Q�����_���?<�Lo���m�95�@����8�o��30ޑ`����-�Ӷ�O1Ne���8^˸��ƭ�����T�"�Ew���߹Pz��q\�É^�/�e�G�7��	O�e��Fg9"�t�ٍ�T���	�;+�8����2�D=z}�\�s��'�&v�|�����7;�zqڏgL�FgU�%��h7�mZI���'�� ɓωyK�1)��ĉ"�sT������RYk���݋���.�L�5�7.���b��h�6����L��� ��H�n����|>�[�[���z2��'ˊ'�!.�9On�@��r���n݋�fAE]�"=1J��ǵ�P`�_�"c+�k�R��4��}��25X
_m�R���f$ˌG], E�%}��YUk�<0�1��;�-B�+���d�`��~�v��@g�E�}C��!�T�w�(fkt�jOm�hx	�|ty�ijYq]َ�]^�A|Z"�(��\_�3d�pq�y��A7�d�G�])��i�E�uu,���v7[o���Ep�%лZ���ZF8Y����aB;䨮�gb+�s�7`�#)�|���t=��zqfΗ���h�N[+�9(Ձ�����m�@&��t�Gq�5Uz: ��7���J+���ywɂ�X�- �sQ� ��J�J�~5Y���n��R���8D5�v�:~��(Q w)��C#;��-�q�StY�Nw�ƫ�uE-I�>�E��%av��~���u?�M�e'�Pna���3���h!¹$��_a�~xS�A8h����f>��:6о��]J��.�D��}����\6g�c��力
ᮮ!-��tGSTc�Hj'���@����.�DXs����ɖ�8R�s��� LA�Ν� o2m����4��E�W)+(sZj�T�_�`p�	��v�V����K�}͠�H��6�miYl�{DbCpZ��e��&s� i� s,��T5j�_�a�*�]�,����B���rq��~T��ޝ��, b8
� |����fM?4 ��rwd�,ϡ�f��bdV�n��9_�qs@���Ժ#�>�g$��W���:�A�:^c�JbpW��\���K`8�s��� Y"��*
�F����9r����dlH�m�Ha��˲����C�(�S �"ĳ�C�w�&����s�����D��C�1A��l{����id�_�W�8j�i���F�~O��(q8��� �����lM��L)��8�X�T鳣�����OE�B&1�B+�Q+�	�g![�Pw1=Av����`e:`s�'��6[�X~"�gɼ*���"$��j�����Ì�:k���E�~��!wx�|vo~p���x
��!R:�Q`l8�^-8ކj�a���w���wS�m 8{J1E����Y���J���2�tc�0\�N�q�%����sŬ�"����I���Z�9ֻ��jmgE�~A�k�U~a	 ���W�>�զ�E��=� Z�a�r?�'�ss���g��.��a.��_A?6��%����/o�*!�6:�0���JjU]eL�q��]T��Z���g,��>9Y�Gf�6�N�-���qпV0��^�'�K�pS#s�},vݶ
L�5z����ZM��i�#B�V�<0���8������7Q��X~	Yg�.��]YFR`�=�8�,�@S�=e�>Z�nʠۧ�Wa�t�FӀS�k'��Iu���#>�/�tLNK��%5���x��Ұ(1l��{A�"5P�'��Є�<��ڈؕ��oA��A&��%g�[��ɞ��l���d���6�m7ޛ&8��T>PARn���Oj��cT>:^���o�.X����y��9��p���"h�ռW�c�Ƃ�<AUU]�;����4;��E�<�KRIݥ�}�qbO-�@k�;�L�DX1Rdͽ����M�gDf���#�Lc{ׯ�@����mp�B��7����i%�y�Wk+��LLU�Z����9�����G��T�w_L�C%E�ץ�*�K� ����f��Z�g]g��U�-ඇ�ce;~�zg?���l:t�dشCUbx�N}z����2�nx��$_��'���"o�"���s�k։�9c�рR
��`�
l�E¹y��dB��jfs��MJ�<��+*��`��D4���,�ϰ"I�j�X��_�K���Hs(n�x�"u�>�2b.߈i�ws��JYb=N$�1"���ݺ�E%0��\�w?0�����(��R<�B��|�+K8�ĵho�X&In�y<Jꤩ�d�LTnL���Z��ޠ]�'����q�)��S��N��|�#;�� g0�r+Z���S>O���IqMq��ɴ)+NZ�^ON�x��~���~]s��� /�u�B���q/8Pȼy�z	�V����J�7,|o����-����9Q������PG�Q]2#�����x��opoa��5�{|8��gq�̾s���K�~�B�;��j_J��#�!Z7� ?#NP��?��T��D��x����f��l=+�>��JU�ᡰ�5܂8� 8�p|���2��9�|@�@�oX ���j+k����B�xW�u��ƽI���Z�zƐ?$ul-3�KA1��Nz�a}�� �U�M�S��
�*e�E��v,�s�<�1��%}��Tԡ�/+_�,d	P�����㱥����e�6�d}��yO'��;�b
4v��J���{�+h�^k9�JdA)_z�3�����s�l턝�[�l�3�#ڐ/��J2i�-��O�H�G�4��}�li��;~]b��������@{�N��b�&S�Z���ߦ(��,P�ɍ�>mGN�`O��t��MTޅ����^���Fb��IN�[�����0����?W<U&֘�Y��^�zzu8 ]��JZ2P5i'QG��,�X?H���Rp�8O�Q�`(�|.�M��:��թ
b������LcF���k���;�_�]���l����+/�~��3�ns\w����	�����BC�b诂/t?%h���n%�i'�q��(��Ͱp�ѯu�-�,��;~P�
a�V��ۮx�0��5:-P�2��A�fT18^�\��}�@}��(�2h#���E��U�VZګ�2�~%z�L�]�H�4��E鲒���5�n_��Q������6�k�r�������w��m(v��n���z?v��^R��OlF���#�k�(_�.]�j˜��Z�ձ�2�p;iPͰ�����z���F��9�V�@YN*:�1�����3�G���k�5d$:u�,8���oI���4��)a��8߿7qK\'��AK~�Cum��^����$(wo��͉ `��Q�ʹN���]K�/�ܨN��b�͆�&3d�������k6�1X�+F���G�E.��>kN�m�\�PCO�թDi��-��H!d���`fѨ�q7+����9Y���M[�K5�&O|���K�G��0�pS�H����f=�[{/���oj�r��ӖP�p�e��Sjլ(��Q��c9�x�[�xƍ��R8�.�n>:D������	���_��c*a��W�;A4p�e���>�Ƚ½)9橱Ӕ��̌�������ѡI�g���?S𐰘�2�XlxV64EB     a46     310�ixu�ʞ���	�d�*�i�p�Ѭ�ci#�8,���V+����1t�-�j�*�Hի�\�׆�ۻ�eB����Mß�0l^���F�A��I&����u�_c_&��LٖfB����Cx�V��ū�t��g"jb�$s�$��X�eO�t|��(��6���=o�C+~2�(��0a�l]�lf�Sw����ƢcAm�����H�`Ǿ�x]}�Ȃ X��Ș_�R��2�9��x"޻���"1��D+��P�w�ߔr�$��c���?�����a�a)�eƁ�ȵ��bc�X�c�f�!Tm�@u�3�_7v���Z��<V�2��Tu�D���6�,#7 K�� ���Yl��2E-�!��۹\U��{� p�vm����>�q/s'&r����&���ϝ_�6�u�B���צT�r���|���He?$�fd1�E;�͵xWxeĪ�&ƨ���c�N�`t�ݦl-�N�2{5[���Ld�Q2�%��I����� ���L�c |1;�a7Q���W/���P�U@Y`��O�VIy&�K<���K ��{���j�M�^�ܶA��8.ܧ����	��m;� x:ٞ��<+ș�|��_�,�w�ht����Ϙ�)7��Kd�Il`�fJG7�.��-5[,�XO��",�x=�]?��S�r������Gz��Q��^���0���MU� �~�e;��Z����1Oh#����E�U[\��ұ��q@O�v�:�u���O��gO���뢩�C�XL�