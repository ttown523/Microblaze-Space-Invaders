XlxV64EB    fa00    2f40����#;{��/E��i用[��g$��!�� ��V����,��sQ�K,|���h+B=CM�����􈈹;�E�qeK6^0	�5�J���������?����@��:�J�㮆��20��Whl�*�����R�l��*l�����
���x��*�q�	������!$n1>�~�?�[gE'����}6�%�j7<�I��	ߘ;��!g���DEr΂�IX��4��Z�}{���J{M���JWC*��t@e�0}�P�sB�ֆ����4�v�]z�o�oJ�m�G f�L2bҋjVp��/��Ol��i�=�[��V���'�f2
|�__�L&���e��c��ir1A[YJ'>�7zfCx�)���%�X��	-�U�\�f����o�˫�eÔ">�@ј�$W9_bt�$��/|�(�7k����X�}Ԭ��n�rE;k���4�����@�}�^����$���rU9t������.ʠ���O�܆�y7�>wd��	�PIo��,��u��S�@{-�k�0&z=e9�˨�٘N��ձ�T��D�]�f��[%����Dg��1�Z{��Y�3�f��� ��ɫ�H�z}���qMa���~�ՙg�VW��@\��U�r%I�}�O�VC�S�(�M`*�Z��a1�Eu�Rzнa���3��j+��Ѳ<��Ղ��/��a���.�խ���S+;K[��@NR����uT��8�X�V�Oe�����sk�xBX[����VΠ��`�E����k9��ݼj�����vB�_��2�r�\�3K�,L+}�s��Gvg236�o�6���`���Nn��i~�y;�q��yx�����%��A �Pȩhq�Y'����x[�(�)*�-0w����w���l5Ĵ�,>wX_3�ƫ��"o5��Y�f�۫�<g$��6�?����Fi*���0�ʻ�1���~�|Qz2���EY�_N�ǌ�Z�Οw�� ^���c�R�$���vKکA8�˂��x����Hq���A�۷�EQ�d�{W �D|˼���� ��p��	����_2z\U��1W���w�.M4'vٖ�I�\k�4��#�!qNϝ���V��
1����S�vazՒ��}ۭA����cx��DW?-��4��ᩡ'z$<�Ɖq�#;f;	��E���WP^�C��>��	GVv���c^g�3�J2�|�Īmj�Uk��d#=�W�I ��N�G�+^6�F	��Y�\�̵3*�aL�]�?gYV��2��`���p-��\�"R��T_���G�l4��U������O
����WQ����Y�������t
]5?YW޹�����)i���~xB{�;�_���>L3�K�˵�M������x�|�}����qc*�%�r1�4���dd8i��l�7�U]�^q�CyF����DQWOS�z��/9�j��.h����|چ��ښ4��D�3��Y��R���b���^�J-���_��g���(s+�k��`qSA���F����|�A#Y�97D��$���\ާ��[���[&oy��n��ج �����|��X ���]��l�u:�(���1�x�}H�D��2vq�fg �b��HǪMk,���#�������WS|@3	�٠:�I��S��<�#$ox�T-���6r���FR�-�L3v ���e����Z;�ީ�=ݩ/��F{�դ:P����nx��9I�uJ%��Q�h��}`aG�R\Ȧ�!ә�5�$�� �Y�t����_Z+bʴBt�`x���O/��;���Jx���c{��sq��)9�U~��J����7�l�b��$r +�1[��'��b|o���-1�'�<�L�"��;�KoM�}��]�����Z�K!,��m`~��Ws�ͱ��h:�|���sA�|2�*�j~�4 �M3��~H��pޓ� ��ޔ<��睥���L-P���8k8N�4����w��wT,Lie���D��B��~��c8�T�G�j>�\��٠g�����ƹH�:	 �[j���q�Q�1��t�a�X&O	9Μ�J��m��Q-�4D<i~"�g&��9��FX���gm����ۚ��i�C���!g	47�(�4�*?�r*&���l�irD�ъ�!���op��|x���܏A�D�x�]�3\���x�֪yբ�B��Dȧ�2K�E�mܘ �W���;��,���Q�^;��NB:{$�B(`�p��2�����wr�;+6$,�*/�8t�O��j
�3!��_U3�,R�����$�O�xc�%���Z\���m^tD���AH?�f��)���O���O�R��~	��D���kyo&4�:&��å�%�<k�1;�Ev'F�ق�����KA�f
�Q�ݷ�M�B��P�~��AjmA�%`��H����g3.�"����ui��rEʏ����|-?��6I�ה&���t3��G�kl��칳�g�dDۖ�Ĺ8t#�棧BS)�HX)��P���z��=�6��?��!lU�v��	��֜p!��N=�%p���$���r�yO@@f�,VJ�d�9xG��cN�S�<�e2,�!=`�0.l�����&���9"��į�O�֟�ڡ>�d�Ɯl�kj�|u��0M��K��N22l^�J�F���{����d%����-�2�p�∊��P�5�f�vc�/©����#ؐ��'�,ތ��t�=��%���'�DIB��u9۾]�'혗6���]�-���m�|�nV�6�I�QB��]��ZB" )��vM��x��b��(?��#�Ȳ(��I���)ޛ���Z/Ǚj�+e�k��W?��9
��|�˟U��#T�{�#��3���fN:�\�.�y��L]�l��We%Nj������+�����sM�I�q �D��/4�]�\jwk�$Y`�v��c��r
�R���D���2��_ Z'F��|4~ȃ���@]�q���S�ز�_��&@�*&���-������7wk�9d"�}���9�Hw�8�f�.꠷?&�?�U��rE7�H���:��Έ7��ȏͪ�lT!�;Ku7m�8Xa����#>fB;m�Ui��6���@�bL�+q0b�ٛ(��D�s�g|��%����*#�D6�}�	�b�F�GM��2{B�qN,������ �+bG�T-^cgW*w�(��0�ӥ�Kff��Ոq􏾍1 s���F��C�,J�OO׬y����7�U��Q�	܈�S���8��������@lԅ\���vuu�����$���5Z�����b/�#+��U�ء>C'lg��S>�.��x#���u�7l�� ��Iaۉ@vߡ��k�s"����ݹdm|$2T֭�x���bN�#-���2��.]���Fs@/������igMݤ�Q_�8�_y녥1��8�[��e�6+<r�
�4gWAN�}�������b�d�?�a�E����Ş(�⋭��=���f��[~���[p%�B�k���M�]�a#�/�)����.k�����c�Y�6�����T��n��x��RG#ecX\j�d�:z���r�z����%mI'6�A,(U޴����^j�XSeX�����L)�R+�G����%1�hKv�Lq���e�`7��TC8M�d:Mx�"oQ��a��]O�SU)]���\���h|3�O����TV��g^�=D|>�ƀ۽�Iݼ�v����7�i&ꘐ�6Ǔ]|�-���)|^3c�H5�5X�_x� ��)"q?�yi���0��+��}����E�a4�^ �mȘ��oکB�C8�|��V6Ō�2�3���ܙh"*��Wߕ��\`0e��T��RP���A,'�i���RWx<�ä�
�1� !����}+NE��K�r(�4n&Q���B>
�r��.���`	�H�*A�U���"�%A�R �9���wj�:����0&.j��{pEb�E�n��ԍVl�ޡp��P�H����B5��6���<��i�S�4�%y5��j�
����b����*dk �GvA�x�QYAep4�6�m�M�*�Qwƙ�,G<L[<�kgiJؕ�
}�vM!�|ρ�-�_�Z�"	��o��UV2�r�Fo> �5�ц��Q��:6�M���V
A��Ρm�<�7��f���(F�	wgŎ؆������Z�y�(�h�B!�1��+l�Gm �8�ڵ*���w�||r��b�̤+�>X�V����zz��n-O��^�9lB���zN���*������~��� ��8�[�H��^q[](q=\|�tfM�V$�����FP����Hְ��"�k�n{tC�@_.����~�&O�bұ$����5]�eg�X zy(�,��7�J�z�!�P�+������2XE���e��D銊H��杹T+T��*ۥ4�B�@��H�8�?��N9?��&F$E�e��C\�����؛ �m��
/�Ï������*���wv��kwE$��Z»t��#W��>~���.f�}��Y`E�� ����.�8W�w�:ו��E�b��ד�s�Go��-�KuU�H��V8�󌊀,���� \����/��	)� O�������=j��sI�O�"��"H.�[��0�J�3x5)e�u;4�ʆŀc=j?�|����)�����g)��m�a����� ��]��/�别������%.�B���#^ǃZ��)�eD��
�I�J�W�
�B�J����ٷ�s�Źg��'�ʄ�x���*���ryq�yJN�MH8\��]a��f伫�͒aH���fj͍���KW!�6�W=�P�����JGq���Z�!{ �!宮r��/�D�8a1�*�p�x�b��Ҟ �H������'��s��e�����H����h��gbT�Rr{h���ű(�	(k��g��u��	����F�Y#����%�T��H�?du����C�+5�s��sh��*K�xk�U0���z�Y�Uk��� ����8�A=���V5=�T�`��"���P��o<�_�-y;��"��v[�78�MϋnQ�)ϭK
�8��A<�Tgv�7���� ��_�9! �y���Ȫ���&Y`���m��䪝�`uI�r�"ta?zV0��)��3*$���:�O���`��P}C֥P�ʀ>i˕�������b������cԜ�h�Q�ve�qQ7���)�5��	���ц?(��2��<��S �^�Uo����b 
�u�1�z�s�2�褳�t�����էY�\I_��#?�t��B�Rm���{3���V�',I���W@��W%��B&ɪ�����*�]���V����S3��A�DS��/�pX��`��D�\�]^�ϝ8�c�����S�9Rb�d�Ƣ5ȸRY޸D��0�����ת_�@�1����R�U�<����n��B��
64�ǚ����VD�^X�z �H��cɋ����?x����߳I�f'i,P�Ne�1�nd���2~Kf8�r�}�ɾ��������;R�ٙ��+�,p0����)��ly����8�FPj�W����#��)/��	!눫��_"�~Շ�Ip]ؼ�ny���,K���g�fM���	K@Ta8����z\Q`�=x��z�ԗ�x"���>&L:�h�, �M������!�)��Bu�f��G�~<��>3�5��va&M�����)�K�B��DF!@͋+����>|��F�o+e�;�z��Rf����L��&�D�"�#��;�3 �$�O]'���e�6�\��#���/PȚF�t�UZ�ۺ�X� ��������!����SR�ڨ��0b��6е)�9?��V�(pm�hy�Q~9+X��p��_A�/ӽ���[�~˷+�xk�:����:�muZb_Fqc�L~�4& d�|�L�Dp�V��6�ݑD���G����*ɶ��c3]�?)�m����>H�^Q���P��6u��:g�ҺAܛ0��M����c�ڮ��wo����F�=M����*o��HV�(���A�4V(L�+FbA�����{������ � C�� p��X�q2?�r[�� �`��"��܀"�����:��;�|i�g%�;2�S�PȒ��݁=��~m�W�"P�P��ktyl�B.�8����V�'��1n5��
�!F��2�d(�@W�$�PD�����֪2��j��P�Ѩb��20�]i�HK�ᫍ�	�קC�)��%v�X�	��[��ڻ;��M����a���=
��V����)��H�v/�m�5�n�����V�l�V�\+M7�J��h�m���k1:���tr΁�2�D�H��G��D9��*G���vW�0#�u����]��{O߳�q���1�F��6���0�1��,yZt�Ħ�J�7Im�~��Fڌ�ü��\�j���l�r�>7�Л��w+�bG2�J.����vy��(k�TmT�^<��Dퟗ��z�d|�p��4����V���:�k-��Y�➳��k���/�����Rq���V[+�f��\
w�
�ۣrƏS ����f��K�Sg�ƺ�6nl�=�-�	t����F�E$=�2[�v��#�&���-�N��n�*Ņ?q�eQ5�����<�k���fq�X��zXe�ReCZ��2�͵<uQw 0\<L�w�T��z9�ԓ�]:J�>��_����[���c�WT�c� �a��aNd��'�i�p���V�Y���,��z�ɷ5�j��?"�Mp:��OI�=Gp˪Ҡ�ˋ��o�����z7���I ��J�g�l\I�:�q���n��E#�ֵ����!n]y�k��JA�C�_�Y���A�^5����_�~U�����|��p�뒊Ry_�8�����8ЦРm������'��z��?ن��;K��yve"��DG�·-�j��;�� &���U�=3G�2��OGJ�.X�A6۞_�!�6��yF��*:��?N>�v�%Iem�?چ���Ox�8sLo2 �i7t��'�����f��/���Ψ�����j�f����A��k�5j1i�R�gY��A�\n�*�"��2��p��rj��`�)�ڳ`���a���f7�2�@�?P��w�������[�Ra���; �|��YQ��$�Ĩ��qO'e
�w��hz<s���~I�٭�%O.����e�d��p;�v��!2�����8�֊��:!�z�vu�f>a��Y����%�z��:��%�}媆���d�v�n#e��YjS����'$��	�:+y$ ��JF��b�uT}-����_��� δ�L��z�n�U͕���T��:^`?=�fu<��c�a�d �_.�v����-�a��n&_5z8�q@x�a#X��cx�$r8���y�K�
�!���b'�����zs9/_�ɘ&���L�뢴B2{i���k�"�Ð,CU�SX#��[�5�L
�t�&�z�9���3��(J�S$�]I����|�9�W�~V����e"ߊV*��f~t�a0䬣��\�0^�ў�M*���iꋿ��<��~����emVv��7N�����It7���"��`M�lb�<_���8Qu4f��KU�((J�z^�&�!��cEU�������:1T �FÁ$T�ZD	;�߮�8��V��%���p�;i�ABSI��kz���-��l�Kja!{
,r�Y4h�(���l�Y+#������x�q}�W�������:y�u؄�?�|�o1"����\�jk�i���p*?��kô�l2�h��7�(~Gb�C���ZLc����.V>w��g��"����j�\�s�Iѥ�`�\�J2Ѣ��^�1ZKޢ��+�c;� )�6���y=���||�>Wl�K=Od�-��Q~񃉰ݏ:��3���,��x{6��8 ��Y���Ƅ����pS���E}�'d��`��x_�A���a�R�x��9���%�8��� �S٬��h�R�ֺ��{��
?����>$}��_����Lj�a���s���V�*�ε�J�U|\U>���%��Y3��B�>���m�c��������Iugm��}E��D�fFe*�ԍzdq��;mP��i��+QI%s�d|0H��	�9��;M/j��������J0��\�i:p���*��D�L�Z�����0��KEL�y��L�jwA�"h�U����ql�?�ɗ)2GP͚����ޜh�n�ำ{u��fv�>��.02��Յ����@/�x�ޡ�(x��Β{Q^|8�q��2MI��~�l���O��h���DAh�b+��Ħ%ѹU_�)N�C�=��8HD�Ǒpa�U����03��oe����U����9 $���hIdO��@6{6��7���/������'���>D�2A2��0`bU�!U�ep/zW�1%�P�ylV�� ꭭�hz��k��kd���Y���W��QF(��I���]�f�z��+�?�&�6��8P�[K����-���'�N�@?�O�B�ࠦ)�a��j����c�-<�ʨ�ے"={͟�4g�jO^��;KC�$NF��?�h�[*��e.m�90{SP�M['q[sE����_�P���0(�4 �zxr�LA�D�uXÈ���zZP��<wC�h���\^�\y~	��CW.^Ʉ���E�״�A��Yw�|�a��w�dD�r�Qv���$&����WY벮&!�e�Zb�YǞ�@3oR�Rg�JzΪ*b�E�z�V�Yo�փD��vz�?�D��(�a�b�F�*���F�Ҍ����z�%�0A�U�k�8E�¤=��B�_Y<E· uDN�Е����9L��:%�l��F�|��q*�V� yVE
R��)<$*?�w�m`��k���(�n;��	#%���Ǩc�e��]qN�Y{�pV`���"�8��
a���9�e��S���i�A0/)�9�W�]�өp�%|L���Η3e��[�l�OB�u��b�� |
pw��țily,i��ssk�qm�-qB|Jfqz����RW䦷�ȯ�2?�W��eMG*��@�������D��������d���@��9��՛�i��#��h녚珶p���GY �~Hs}<n�ZN ǋu�IV�v#+��w�w�)?��+�F� �S�i�, S�~;"��+����S��7ÉaE�ǲ=h�݅�u)d��0�?�dql��a6����7��0Yf�<laq�2ʪ& ����4W˿:�z~�v����Lٝ�>q+��i�u���QJJV(��o5ku]d4�Ct�	���v��I���	%~�30�j����"������?}�h/EƆ�:�:�s� &�O�.=��.v��={�GL�������ez������$�`���-{gvd�J��+�[P�=���wB4�t��p_������D�AX�4��)ǈQ���G�-�-6n�[Z2�uYT|��(�C	����9���59R�oȉI�f�xd��9���:�Pq�t'�F�\���(�F���A�Mq��0��R5�ꆰ,�ѹ��/��v`vTRśẌ́!P�{p�,�`#�!�*o��"?��4�\!C*�_�c��VXkv�'�����t���0=�%Ͳ5ހ�	 x;*j<��r' *m7*��>sM��&�C\�#�@=�I�	�e�2��?��f
�����GMX�Z�ZP�@��-|n&���b)���4�u�cR06P���y�]�0���St�u�� 9i̾�}�+]c��^���g>�ds���.ͫ�M�v�$��S;7��Q��P���l���	�!)=��c¨O��I��.+���T����� im�h���P�YG���
9�BwgE2�1�Ȋ�T7F )Z��n\oӖu2�n�~{yK����<iY�ߨ�̰
F#N4.��x�\	 ����Cj����Ñ�@׸�E�$��Vh�9CX�-z�dв���@I��֏Ā�e�c��{�m��qd-,�I~�*���B{��o��[_��!R�����E�8K�}�59�>oj���|�U3O͹��<�͎��0���s�~9�8��K�zS�ĵMr�e!�"��iMJ婇��`��Q�7�ة_K�����~�����C��j��e.��1w����3JfZ�3fʘԪ���������b.��' .f�A�e��<*e7��H�@:���T�?u�BL��X��NapCӆ�05�t�f���lQr�1!r�"���UL<u�\cvD�Q�~�P<���㋰���@1��:�yn෠pw��|gF�MJm㤕��?ϥ�ųt|�׎&�9��s�C��	%t����N.`�+>��Ux����d��:j
�L2�/^9�@A(��?Ƈ�'����,�����CH�]bE��AdF�{��57H��hY7؝��$���>�\��ͮ��hݣ�D��Ʀ�c�E�@�U��dʚ#�{B��R(̒��̀b���}Yp�D#���'���� x��N*�%0�{^�qˉ�p���~>J���uƉfy�3��7�U���儂��mDБ >�l�>Ʌo�Z��-N��A<ZY��Y"A�A��M֕6P��e��4�ik�G(���!#5[\R:{OB��y{{Sr�U8�8Q�&|>�ٍ�4�n�Kv���(ڐD��.��ѯ��e߇cA�Z����yPֱ�-˒PP]IrnYa\��G�\.�-W\����/�_�
�e�D��tqR���?A��/ʥ7�b8H���[ƀĎ7��$|D-k9o�.��8��Mʼ��P�U�3Z?H����\o�=�$��Dq�F>�?a�����w���D���i�ђc3�µU'lN���1�a�u"._mj���7��K�E�߀�3��G��K�\%n7u�C��2�~����m8-�BV�ř���$���e���:=�@t�b�E� &���+�����n�$}�~�ȸ4؀�խ<uYeF��~��žt�q�h�8	j�q�-�0���-@ ,R��r��==�����~&�9�/���uJM����w»� �� ���F�������{���z���>��.��c�K���	#7'՟Z�I�x�I&FJ�7v��"'?
j�B��ˆ�?,9?y	��mo�yi�*lL�>�J���~8e�U�ل=�a�h��V�e��*��J�B��V[�a�DK�-jI�w>br��S�Ǵ G���cӈF�n+���_P��H#�X�Ē��dCƋ󙛮�)����#؂�_Ӕ��+�9�#��r$�Zrvޣ��z\�Oth�sr�k�"�#.nb��$)vG��������\�+�0����ʀG:�O��Ĕs��^8l�S�z��k����0K|~>�c�?u�[RW�X<�������f-)f�1nW��鮂9��y�'ж������dX�{Q�g�������1h�\4����3CӃG�>���t�ۛ���SY�g@�$�y�j_�N��Kg
�-��l	�1Kl��`��7�ì���\�O��R�Y�V��f�	�Br�٥�ˣ&�\O�+v�q�j�#��͚�`X�`�D�g)\Ng�S��˓�ݫ	_�L���-q�jڞ��w���p�)HK9ʕӳՖ6�}"�EvV����9ϡ�[������c���u_��a�Ï���x����?lK�MM2	m�=�LO�����K8�=���i!W
֧�kW���Ao�������ZL����xE�p���MM�����kj�BpO�U8��\�Qs*���P9�P�!���;-:�o�K�_'
+��oo'lW�&g�+��]��a1����| ��3*O%�_[8�rx%����a�"�cZ�[k>Mdmo��e��ټ���1vFa��1�'XlxV64EB    a643    1be0sXap~�9�e�)��2�K��f�Q5�&z����Ѭ���d��,P�/�����!���5�]�C��7}%��G�[G�1wt�b'O�a��Y@��)枦b���W�+:�����Db����ŗ��*:+�:y�^��6�<���qu����ş�s�Y5����~��ȭ;&���r;Oط��X�:�O�W����"����}�{6Y����:D��l��z��;(Cg���e>�"U�z� g!�MfPw�:��t���� L����R�o�*OkW������6�?V�����8�yNy��R��'���1=�k~{K#F����z���� a�I�pM��KV[�:x��d�>@��qrl>rg�hN��5At��?^�Nh9�{�>�h��6蔳`,R�h����w�2��>�Ez�	T��aN$>C MnA(97Ni�X��}e�w�E~���,q3���VU_P�`._�k����3���ك��X3���k�4���� [=nD������d�].�Չ{���܁�O�x�1,ݳ�3�j��Ѽ������
L��y�j���PJ�����; e{�b��B���,�¥������'�FB�e��?om.�J�u��<���i>�/�*|���'K��p�\�?�CY�wD-�kh9�o+�7�z��S���7,���E5?H4��g��L;T˜�����KHB�nt=3[�O�<`fyEQ���I"�jzZ/�2b�	�"�j�� ��4�D�D�$�-�R�=0��F����@݇\r�p���ݝ�9כ�e�q^;N0�$��>C,�Q��@�%����#�߻��+����
ޤg9R
rZԡS�pOLdڊ���5R�b�ЗZ_E�nB����(�Q�G��W�di�DM�
��枭b�����h�j���8�Jȁ���Z@�M�krI�*;�sA1�d������*JE%�<?�#���xu�ʊ�_��� ߆����V{TP�~-�Lޕ���/�bFJV�����#*hYY#ap����ک	������D_�x3'��~#���)n�8�S�3�융چ���2�Tu�g�3�+�/W�|��\��`pý�%�_���.�Ep��}U=�GӅl+Ī��4�4qw����U7g/�D8����0!U���j��۶��g|MM���<��P�uoz��0�I��K��h��PI |�����x9�k�E@	�v�ӆ� <�ZY�[�iiX؜�+hQ#��{�mkՠ��;gޖ�c�Ţl��?Q���(��ӰӕK-28w���T��S�?7�}>|;�N�o�#�XKo���u:܎�>���t��p_�W��Yʿ D�+����HI�V�%���ݡ4c�;� ����+�sÑ��(1$b���i�a._֎�%�RxD�Ze@{g�tI��ݴmy�b&%k�_	���#��#��4U�pd��Ч:a�#&��pCJ�}Ǉ]M��*�b�ya�R�n���&�z��F�>Tn�坦�={9s`M� d�����pOC	O�@Wm՝�@|���f
�iG���Q��q 81ۄJ��thpZ�샿��?�a:�D1�@��S��澘_�T<�/����D�z7ɰ����M�P i���� E���ϛ�~՘�KT�E��R��q1/�z��4�D_�O�h�o#2,i�� ���
��l|-'+W+�ąιm�4nS��>.;��+�����S���_�Z�s16��&J0�Tӛ魬���$�E�����,[�K˛�,�{�8�1FNB�҉�YL.è�x���0�3-I�6 1��J�t1p��¨jc��컐�:Z6���_S˃�A�F�s�ES�C�r�:诸���X��	Y��)_,��E�r�MJY��r��{�HGl\��k����L�(���V�[ML1����y�x	J�j ���(�N��]�ׄʿ�����Rƣ��,�ݔk�4�*�}'���((�Ls����B>1	��oB��DG�!d����3�E�dB�`���zzG� ��-L���z��R&��_���Uk��0��
S�ǻ{x_~o��̎�/�ہ��:#����� �3y&%�?�'c��@�fS��R��cl�Yq3��:^	Z�K��
Y��M:�2,I�^ф�N�U�c�Sd��C����S0,��1z:�~VV������m�2�+T&F�sV,������o(�(.YES����P�&U�s��r5!�zI������+�
�/�3X��Z%Κ�2� ������<���`�Q|���^���qBzcr��9�&NY<��8�����їڃs�{�U$��'�à�?e|��Wp�hg|�/�ܲ6/��=��P�M�'(-Ўd����|���iziG6,S�E=��>�̙l��zmό��̷+�֪���Ǟ�\�YZ�K���LkϹ�B���T ����9�}�=��Gr��,�O8,�:\hlU�����Ӵ��;���ѷФOt�H�H�:��r�I7��ac�W�}�mx���>����x9T4qaowoFM@<�Ȧ�-\O����K;�,huO��į'^אs��6�8�a�o�,���,+x����,�������CR=4������*�wC1�Dj�М<���_1+��ӤT�b=���5KH��K�w�@��0{p?0t)�lc$gM)�z%`��a���6�����Պщ��Y\��0�?hQ��m��設8��)[8��p�6�3Z��=\y�a0Dk[k�j嗾6�c���2=�+����Ř��P@#gS��÷�Z_YlN&f�]G5�80�i�%E*TuɓW�ͷ��p��H��R[M�,3��%,<�yl]|�%�^��'W�+�ƣ=p�0�!l����5��84����{0q@�ӥ����A�"0���j˳�>�؍8�������X��vi3��W�"
�]Gq�u��$ x�3u��i��0FP�xԁ���T���[K����=rC���l=2�o�+n�9_��dE�,�S��4,���?��i���c��(3������5\{����>G��"$Rs��B���=��.��}�w5�����:�O<q����:b,Z+���������a��#���bu8e#w�?|>(���u�&(l��KvSW��($�v6=Lq�)̲g�C��Q�7Ѱ��v^?HH?-�{�?b��-�����?���}?����,�%VR��#T�H=��R�=��W.O��	J�4�<*D�E��O['Đ���gM�E�>��=�EN��[m�V��X���U�����zo$�&��,�%x�)��YT�fk�\3L[����=1�-���e}JG6��!+3T��\�'5��t}��]oc�f1�U�ڑP��*��[\W��l����զ�� !��v���R��`7�M�P�<��SHl2�1鼻��՞A2DM}�w`�3�֋�p���5
 AN\=�eiE�jR��W;�WoH�,�||���\��+g4����ǜd�ޚ�����4���
ܱ�����P�O&�S��d�k�d)�����,G�JNӯ~ue�B
��ݠX�p9�t�l���&���}���k��ʎ	y�̄)\T~�(b�?*ٛ�Ѯ�& �t�;�ΐui^8��ޚKf3�n\�hi�/ۨ		וO� �@�7Y4�|<[����ME J�s��)q��IN7>O�Ӳ
��-s�����[��o��	y���Vt]ޢ3×��[s��7�/|a�+l3V$��+8_��3#W���LB����/!.,���~��b�����8�Cڼg��K��wf���@��- $F;M�R�=V����n��1��Y�F���4WI��>��!�é�q�(��)�7 ��F�Xv�ϋ�ab��9�������Z�3K�0�?ey6���g���w�@�T��_�4Íh!0����[�^��3bm�hGK���jʴw�$I��%�l����`i㛧᪩S»'�k�WG�|�k��'Ժ]mm��IPO{< 1���$_�c7�,n��j&�~/������f���;�>�hdr�����p�[D�
m�ޭ�{z�kk����&�3X\t� ܴ+]j��!���V��5�tx�;
�"�L���}��.۴�_�O[����9�is��b6;�|����z� �͐���F�a8D�-������ �n3pB9Z�
��g�d
�B�J]�&:b�]$��b������R��2��ys�疝�4J5m�k�#�
CKԃk�dH�A{q��vM��[v��Џ��2`�:�10���էc�*o���(���#�K3Sp]؃�J/��Jx\����bb�DR��y��>��3�&����/d�ҘA�T4G�g�%�^צ��v֐38��D�&�4�KI��/�!SC���*҈�j0��n�c���E��.xe�#Ի��
н1��(�<s0�".�{ia�FAqؽށ>+�����[H��E��E�<	�7�dj���D+�#�r���e�^���5�;��ފҠ�<2����� ��f�t+��ޣ��Z��ӫ�EἬ=�Ws�6|�C�Ǿ�ڤ�.OX�e�{���J�=��C��Ȱ{f�W�!��4gkA&F����� S��&�x��xȍߤ W�4�*���V>�bR�Z��²+���QN}����'c�{��Rqp6O9r�F����C��5��f�8TA�����jޮRi� A�B�����t�)���g��4H~��ߣ~��3��|ʨz��1���]�m�N^�%CI�R��s*O�$e|�e���/Y��m-�_?����T��	N1�7[��Vp�1&S'�����#�IdY����&�c�i��!�d�tfǧ9�(Jv-b���r~Q�86_e<�Fo�!K�m��r�%)o��W)�x��,��z��P����W��Z��+RJ��TP�0맜��j�:��[�JDs̗q����WT�_E��ϔ�Y_�@2V������o �'�d�1���/۞�6�	��!���A;��cԗ����k��Dj�p�ΐ����XJ�ڰ��B�#?��^T�)+fu[IC�B��x�)�O���%;��"�Ǉ�>]Shr����_��ڂ�S�[0Y*Rh���NnX���!B^���h壜!��<�:JkP��ID�v2Os?E$ϞdQ)q����Wx�q���h��$uqqK� ����Qz�Fn%��/�A%����w�y���z�[o����yi8�^���#Z_���lM�rM5>�O�)<��D`�
͜�/�A�:_�DYN	PC�&ovQ��b�+Jb�]ԏ�f��y��M�Y�g�Z1�K!u�p�B��27ߪ=b*��w�����]���~��2�9����4c�"�eZ.1�_a��S��.�^��k������u/��R�PD��D���T����b���!{����i�m6F]ۻ�hujN~��r*קW��r����9�?���e#��J"_c��F�'�b#��ƫ,Kith�rS�v��F�s�����t�x�m�/��mM:�ڿ6G���ADI��i��RǦ �t�c��8�#"�5�M����nG'�,\�'$��]��{H�Fg�O�h�rkX�ty�c���/ek�t�g����	���!���J^_;���HI�{��]}���!A��b&W��hzesv%��k�$베P�H[�$���)F�D���:��1Î�[�,�4�p��kU�`X�+��I �o���zdY+��fn������B�r�6�:�x�=�2���lWo��?�m�w譱������$N�[��D��^L�o�o���pO��ܫ�]�t�u Hy��Q��s����$�w2�%]L�!H�v}k�%�n0_mR��wgkK �A�e���2�zn���.��ĄĜ@�4�w�$��@��v�H��#�zr��K'�VWVԸ��+y�Sn�G��A3��`E6Ы�p�_���N����5۔'̋���r�)m��u?���H)_l�ћ�h�N`qx�WYRsZ�3�(NĐpN
���x{MR�=�p�5-��N�"2!�}�����0��a[[66Rg:T���8�Վr�����5�ȉ�B#X��e�;e�О�Q��.�ͮ�!6�鱖R�S����	�wT�~�p���)��3���D߰F���9����V����O���%��oB�6kZa���q'�(e+:�F/L��F"z��sx���}��mY��x�� 0 (0A�> ���}̛�爮I����A �;��Gc�<�G�qΟ�/D��5��o$2�væ~�\#�@�61�h��`��(*��T��N���ʽ�O/����_C���
��t_��ÛZ��� ��jg�aV��H��&�C�����6��s�@����2����`�Z�"�NӮ�]�ĵPYQ�Bi��Ah�NE;��7nׯ���՟X��^O��u%��}_����kZ�`g��~��Qwgq@%�M�nKǵ�*#����X��(���ٮ*�����6�@�U�O�-�P	n��k@g+�yU�e+>��Cc�|y.B\jr7cP�vt��1t	]	J\Hy�[@?xA=K`_�R��``�&%<2��BWN8{I�NZw�fQkd�ⶕ�I����n�H�ͼS�ව"�_I{eu�6�:��΂�VM�0�ط�*����b���Ӏ^{K�\}�0 ��f~���������V���Η̒��=�W5.�7��D>HI1��-���x�'���RHY�AK�R��?Y\ �z�_tt�9;�{��.�#D�Z/�S��2gIo��r�da�},
�,42���dͬYqV�-���U�b3d��D������37Vk�X��K��>s�m��G<�cb��;�}i��N��v���崎XFq�R��ٹUtaf>���sCPl~��D(������j^���Y���=�x56��?f6{�v���s�>�hY@�| �̓5&&<&m;���^:$c���+oq_��1|�5@->~mYP�5��Dx����x�(�+����Z�