XlxV64EB    fa00    2ed0�#��Ҩ�Rյ7��;�����(�`l�s�.>t5�&Q�2� q�$N� r�P�A����	e�*���S�{�MO���?��/�t��^�\}�%��C�u�#t��>�GDR1�b5[B磧�$>L��*%>��N��W}~wp	���o��>{*ɴt/6��y}�^Vl�6�N\(����{�'񹽾|X��~�c
�ೠ?R�Z٢����r�B:�*�m,g%SZG]�k�h����+��P��(���y����n��䛋T#[:_�?�ɻ��O��	1rJ�ɨ��^�mq�P&�3.�	 ���D�Ϟ���<O�r�_�!p.�%�<��J�,,m�C���HCJa8��-M��h��B������eI E������C�6�m�3ZH�"�9J�z*�Q��H�gw��5�m/�������,�_�B�$�D�e')o�iȋ��P����5�+̏J�bF�` ��=���O�"�L 3y�b2IP�o�!7uR�G��k�������w�\����"6)ɴ4�7�+��$��R-���Ug��@��S=&����"v��@�:� ��C������/��{ƿD�(�L0P��ۿ3lK�Slil�Kh*���x�$�3虎U����b�}լ��؋��I�����0~���Kj������k���<QپSQ��J�C<0K�Y��q�@*n�����R`C���4�I����HV����ϙ�Z�O84���ؘ���8�RHb�t5�Jؼ��ţSp@q��Z�����I���d�%�����g������|v.=�p���{*X�&@�!�$A���(�&�X�
�O�K�ɇM�ǩ�2��Nbc,dvI��G�e��B��� ��Zu5�@[��8���2��A��3�K��Ǘ9gvE�vqU�����w��3��.�{Oc�!д�~sX���?��<Q�Hq��P��vjV��mԹ���%�I���#=O��{�5��J�Un�]c���5���Y����C%���3*m1�h�rd�(?�k�i3�+�>��Vs��%�H�ß����v��QHv��� H��Q[��j���no�ٺ!	h2J�χڬ�eЊ���Ƌ�̯! Ե�t}�$�Q#�9E9��]�A��v���Z�k,�c��:��ʴV��@�%G�e��J��R%F` =��еn��3��a�ƚ�g��R�K�����2����)�]����n��K�J���l�x�k;��-�˯k���-�Nq��<�3�S��B��L�l�I���}�P*$b���+�j+�������GBJ�W�UU��A����؅��?�MYnXw�	/p��G졵;X���*���E�Q�M�u~�����,���s��h�u���hn;Ĥ��?����ϟb��[�s`�+q�*�Ȥ%��H|��C�;c,B�|z�x�:8$%���~23ݎ �%�˲�k�C�}�E9�r�*��Ld������n�'��$x&#f��=f�2�k#	���ڔ)3� �Ĉ<3�{�Q{V9�lsQJ��.UǪۉa	�����b�*ϫ�"�c,>��y�O��/A�m�T��֔��+t��C�&~6o0/�jp�o�|��ha�I��f���n�(Z�H@e�$��mV�Ȱ@)I��߃=��3p�m��7��4ף��	q���u݄����E	����^Յ�	6^�� �X���8�[��WuvXgQ"�A����$dA,ҩ4=���Fxa��$��:oOJo]?g$��@���KL|�.�b�؇R��嗡��~�`�/���V�eD��⽼|��Ƥ�X�.4�mB!f��U+h����N��'I��`K�[��K�h��M�@��x��0e-�Y�[n�\��I�+
�������P�'��Q �6��i;��)VH�+ފ��Q�6����E�_���"W�GZK� �;HGط�e�L�jU���b@mW��&ͨ���2��%��Kɿ���4eH�_v���ԑ�V4WEb�Z�Z��{���POם����:#���P��� �^3cQܑW�+U/v��F|~3! �W��u�fĝJ�'d0Q�zL���M&6�g��h�C|u��-�ܗ�D�a�W���U߳Y�7�-]3���C�����&G^`�E��3�]L1���������F���:&}BG��C���"��WNě+���ju� `����"X|���y�ep�������Jz��c瑅�Wtf(�V��M����V�|���!K��t.@~h��-XϦ�3p�����5��W��*�"^�>ЀR`;������>N�G��דXᙄ�n4����ݫd2#| 3�Эc	��lJ=��A�՘�ұ!@��R.�ރ2"G�K�4�ڇ�F�t���Z/h�H1��)�9�=˨��?����{�n����)�js��0���§��~��V.RC�U�?���5�Q��ڨ�HEb�������q,u9��4����#�$i�l�U�=�ՔB����֪���B+,c9W�X\����z�T�=4�L`=��X6�!�R�#����G���0:2~E����mkAB| ƠC](��)^^|Us�%	�#�6�{�-��-�)�8�W��\+���[�X{��ڵ9P�U�Xjq�j]:�{V.಻zc2���������_B��
�g���P���R��g���'�̡ �y[@�W�5���{X
�Pb�`&�0c�xlv�ӑ�V ����r���8z�����Ǧ����(�)�����C{-�&�&w����Q���2C�}�h�4�6-r�)��Pds��Qa�f�I���j�Y���D�"~��a�B�>t_�7?j5�t��B�����N�=��G��1�Ǔ�`�$�<=�wb+�z͑�����V����V��p�OK���������%��8�������3�[���X��㜡�lRsߕ�{��b!MԎ����ئ��Aԋ�{�����K N��d3���>�9Z�H�Ӗe�,H��Jv���MJ6����4?��7ڊi�v�td*Bx8�{j�_.j���E��*G| �b;'��i��3�Y�\fDcO�	����6 �Y�"����yն먛�H��ЖK��D�x�r�VVLHn��o��'�B빒�9��~&��Hĵu��Yi����f��ç�l�h��Q%ndUY��Nc�֝P��LB&<�ᄊ���I���B�X��t���W���\�mA��8�}5��z=��P�̴����<^���0Stv�d�?�bBR ��D��<9ɭ ��ri�`|��S7$��g���
�l;��}H��n��ϲ���moXLr!�g�i<4�Y���8�Lc��M�i��hͽ�T���L'�,��-a����$M�6v8����®��L�hA�hDa_�s��x����{?��_?�z7����"7�������=�"���-�my�"� 1�#��qe��p��s"��W"9k8s�%2XQ�d]f~E��_,D�4��D�B��g��부��e����K��<�*6$h?h�X�h�s�֞�
ʛ��~X��-PJ����v�>$)A�������2���+y5G(� �����nAхe-'�TZ��a�߻����-�L���Ei�J;���O6��ea �g�5o[Q8D��
�o�������/,X��Qgͼr��'�y���'J14����f��Y����5��Oq�8{��"�C/����s����g�?�^�[��J�;<8��l ۼw�I��q�^��p�ԇ���d��{y��q��ǰ,AX��q����6Q
f�=�=^J���"��;^�R�(� �}�uSRC�-������D��������R:��+PKe�н;�����?&�� ����랡��	:���դn�֧0DY��O!� �V��D�'x/���ͶE)B]d��Q�9|���0�0�o�%����)U�r���Gឧ�M�҈�w�AL��W�kŴ}�@�eZ[�)7(�X�W���1�/e�v08��*��YC�aT.:����uՂ�����0�iXR@�E�K8�d%�O~O���JA�̒��_/�%�b��z�˙���T>;��}k������Z�|�9錚��/�Vzæ}����TV��N���{qV�~��*z���R��\XBPS��p"K�_�!�u��m�	_E�x��O��� �,E/MC�z`ͨD��a,@����)d�9ъ��KQJN.�9�غ	d,5��s"/���o}���L���\�[	��6G�!	�M���L�Ln�E��n�l$�p����aӌ{a̳:j�O�F�i�Ё�`�V�9�=I0�=��X��c�<�Cg�=��a��N��4�A�-����U#�%��f����z��Lb���Z�sl�j�Ͳ�*b��X;�W�S���$���-b�-HAKY=���!�O�3c���ٖH�|�
�ҧ�����R�����Ї���q�2�.h���m�N&1c�
�b�p�cn�>���L�`:�3�����w�<|u[�Q��x���SP�Z���Js �� �W��L'B�А��K�N޳#8N�<;�� �M%2V�C�ڇ����_۪F!����/EeQ�1o��(�?�ى�$��c�S�/��&��'jŒΪ�<�H�[q��%	��V�Cn ?��ۓ�X��6��u`e��%?�w�y��>�=L�p����Aەq��;�Hwa�̼"�ڀ�+.�.*�Lx�KBp`�%���5@�._�!Z��S��23Ye���.��5�⎴/��O��X���ָ^ *c|��nւ=In*�-����E�_�-m.��1CDq�h%�Q�pA� *�6J}FXa�f�SYGZ�\�n�g}�<{~I�cf1�%�V�%�h�Qw�+N6h��;�`���2�ty�SrQG��L�Οiq+ran��Y��׭��?�k�P�K�`q�p ���	�4�J#���֪��!��)'3ƛc�˒z�1���+s�ⴹ�4��̪�e�芹�B�aW�J��a�%<$��?�33���B,��;��+��`Ű&���v8D��ȅ!�]���򲨏wb��q����W����e�dG�+d���G�C`�P�<<4����ܵ�
0���^YU�F��n�	�A�֣-x�qF�R���z
7';҇�_Q,�%"��Dmπs��up��v��e�Ƣ8J|��Qmk']=u_x��t�X=��`�@�PK��I1%���夳ք�L�po�:�=�ͳ�Y*C.K�9<ґ��oK��T�V��&G�h���H[͉����%�,��W0�a��һ�nd�[��sH�2�B�`�k !s�!,7�!���Mv}��L$xmY0#��ؙ��~�%׹�+``K0�Y���fB�""I�3��nF%]��ı����\��NQ۽%q�-�׷�E���E�ۯ�+����x�j27;4�Q�jT�C3Y���w3�F#��]�-�E̛�J��'enhk��}�W��W����/-`<ھ�?;������M�S��ՐP]��4��g�%���+��M.�1< *�j9o�����7�r�YTӬO�N	���>�7{�=�k�`W'6�A}�1�>�3�O����f
n� ��N����a�YE~dm�zW�eڷdZtD/�E����R\F�KxN�w����0O>�7����O#�r��{+\F��*W� 
|;��7��p�B��i����= ���4q�Tt:B�T��|X�9�����&S�O�r�|��[�?t.��O;��|e)�F�����8�AȪ��T:u�n�y���v�^?keY�<,L3(�<tr4����J{]b�k:�& �DF1^ "|V!���^|�h����%�V���y��z�����V]�ّ�'"D�Ҷ�\�G�'m�l�H��jb�&�	�R^����`����ɜ2Յ�Qy�8�>w�;���1�*u_>0�'�y^�]�V[��g^�|�8���(U����5G|ϾGv���u�NSi�J���EȬ�m@�Da��e3���j����_\.��dk*�J�G�>"
b�eq�˩��n1{U�ǅ��,���'[�^tܽވa�cX0�s#���z�%��'T�dN�y��k�s*�:e#����<B����K�o΅2�f6z���޵;��R��N�\�:�]�瘂͵|\.s���f�/��?^:�F�	�J���������`Z�r�1�¹��Tq�9�Cmk'�%��>�,�	U�VI'F��H����o�i,_�X$�����x7������7�d�@Oş�f�,�(O1�m3@��q'�K��grA���(I����[˂6^�Q˼]3iX�������4�F4�^�1
��1�Nm�O�~g:��W.p��8�,�l��"17_��˕�/��Lb_�� �T��<�Y{��<��S��MEI���V�Z��:9NKpi�)�yI���¾�������堶^�e��Ja�V���4����.R�o�&dX�s�S|�0�B��1ԅa�6���\���C���)}UDqkő��>x`��c۲(�f��`-Rdq60�mcc��kk4�6o�� �a�;��O�^'ѿ�Yd-=�ZĐ2�M>�-i�J����3�t�R�+�A's� ��Y��+i	�4@��ORL����
hA�z!W�pz�+�w�`D�Ͷ�Q�a2 ���&v��L/�'�Տ���g�pi�����%P�o��+	"^KL�/I*߫��_h;�w��3t���HQ^C����L���L>��ķ��]j)B���H�~�AߣB�XF��V�!����qY�C����Th�i,�1 ��,D�ɟ���O;|����6�g%��U�Sf.�_T�v>P'Ʊ�� �]^�:�h�2�j�Y,Ht����0=f��J��+�'���,#xDY�Ɖt����j4�ofͨ��JiǊ�{.��'�� ���� �n�R�Ն�r�g����� �L����NM���	߸�`%����u����7j��7��~�<��P �9ή�	^f)�Z�]I����w H��iބ=�H�:��|X��5�o�ã: gzi�E ���jN������-cV��t[-�\��bd���ũ��ͤ��z]�+⋈�r��p�,5ф甄�9l�e�p��>�rry#I��mFy*rcyó�fcx�c1�o؁��1A�	�8$?�Ӿ���Z�S�5F`�r;��Y�������o>�t=l�֖!����r��䴍b�c�Ofl;�=��:z������W��f�ʪ<?�oi��8V��\�D����ZX�@�6�JN��@k�3 ��+��b��ު~h��S��=&'K�������G��j.9�wA}P�R��e�[�提�R�D����8?�p��n��bW�����؅V}Hܙ��B2�K�o�ʽPz�o����"�<W�}���j*�]kU\�8����t�G;�6!�0��c�y�V�^�ɪ��t�ͳ�tx�1`U�}��{�@v*",�dA�|���C���XMdX�2 ���������P]|H��^7F���$� �sd���kD�h&򚥐�G~�N�{Ƹɜ88�y��d����ɼ\Fu�*7:z=��,C�$ﭽ6i\��%;�y��J)w��Pʁ��D�Z�����w��A��6��8�<��� �����sO@�f9W�~�g�}oB�*�"��F�� 3����gJό�(Gvh�o=�rF���Pj-�M��<�_x�% :�3�i��{
V�_Ж�"�f
�eR��A�F/��#u�
nv�T+��w��:���e���pf�Ys侊��>Q������_v���g6�`� (�B�� >�H`Ǔ��M[(Mq�7?*3r��/��Ʃ�y�F޳Ji�E-�D
٩�����"��Z tڻ�-��W��/m�dwo�WzaP8��T.Wr��d��.g,�� ��bƋ>���~T�"ƠiXެ����zA��_���z�7?��޺@0�s��&�)�J�pj�?T��̈́4v���afJ�quP�k��-�:5y�	B\Ch/��JB:|0�&J?�~Kr��a�>�p�V�Hp�����<N��?L N:vL��lÿ����������Z��%�2�����Z\��`���e�'$�ݲ>崾z6Cn �4��>nn�L��2qT�L�Cݦ�Sf��u%�Z��B���S���\ b?n#	p	��ݥ] �,��	v��a+��D�-xd�_�Ic��E�_��҈R�<�du罘����;�n��Ջ׌�fg�l��>���`���Z���WϿ����G�ÈE%�_�����dyrս^�;�X��8I�d��!D4Anx(��߫KP[�H�Pxm���n�o;�ᵢ�*�9�c��q>�j��&�?x��Ī�Tx�	ı���/����M\Y�*xcn��O�* �>"a�T͛���7��e��w��#���~JYA5��R����V���,<�`L���|7�ߧƃ`|W��H�π_�d+IT�/:����c`���oc�������K!�1ۃ4��ХQ��ū��b�O�k#k[��v$f"�;7�=4�5��3	�/�%*I���}b��������*Y?����v�)h�p7ˢ�1.1�@W^������O�^P-6�%~�-��IHmQ=ubL%��ж&�,���|�O�<���4�~���=©)�7%�Й2N�F^�jS�ׁ�59����oT�Q� ���ݛ-�����O6�d\��ª�z���r�\�L�Iz
�y+׆��}��3W�!�H��M\��7��<Kߋj��W
�dȔ��O1�xv5yi�ƽ�C���z����=��A`j�NVQc���LEM����(۽'W��^�����c� � 0���FG�l�o^+�:RE�(�[
7]���xWdnP�-��!P7n2��~N͏b섙��bL�"E��G9H\
Dbޜ�����Fq,�� �z��^(�����{��M�R.���4��t��~��8�Z
Pm�7��sA��P�Y*`���K �.Y���x~�7�]Y���� /���]��iYZ�]Aw��6��H:�rT��}�˙+�]=tN$�'���u�$�).Ys䏚^���G�0��ڻ*��m�@Q���}��F��rA�Wb_Ϻz>��_죂��Ds�$}�,x��U4��z���T� h�	�-EA�ي0�OU����i7��"/NO���,f�_qA}�Ų��,� f�:vy���.kх��t�W.n�D⌅�������j�Od�@���/l�	��VLB6	:72"6	Z�(���������s#�mbhK��u	4ʉ��KHJ K|��j�\��d@��֓����r��@`5Z-�Or���8F�Z�1b��쐿o���Gaq6�0�=n����Pph�'�A�$4��mZ�b���K�X�i�I-�U�gf?����UV"7�����0E�E(�T��&�4�ʡ�ل"vǾ��f��39R5��ջr�J�~A�Q"�t0��P��le�$8��k�Jem��nw��:�H�/~5��@"GF��vL�[ou@,w��jSb�;����f+@>ơ9���^� �L���8ZO�,�?�IB�r�\�^"�~�XpC�f��t�W@��Pߌ\
ߍ�ذa#���s��
�Uq��oF�eƒ�7������t�L��?�,��AM������}�����Qb����*��^��ue�K3Hn&�*r�zz�z�"��(�v��R l`D=	`#�t��� �!���F����I3lQ�������}*kJ#�ؓ
ˊ�(�/�i�m�V5��$w���Go���z���@�=�#��{�QZ��R�W�7e�w�H��!���F,Q��ѓ^f�,BE�����\p�|C�lRã�~�1+O�6]��"��,�0�ݰe5A;>�bXp����C+�;�l�xm��ދ��G����>�=��Nрe��\^��C53?�'����a#.Y��p�m3T�̑2�5�����ժ��XW�(�`ċ�r�.��ÁL�G�)�����x����n��}�w�6?
�4�d���v��Ԣ�h6y���W��?hg-��y�AUC��s���υ�i�qi��s�
A�R������b?�Z��n8N�m�Է@u؅4���eE�<�̉3پnν���K$���]�W�!5bo����������9�"������l� p��ѝ�?j�O�Ƙ4��.5w��|����*�"�k�PEO�Dx���@f{ZB��Xj[�lRVq���RA8��a�$��*��e&!���l�kcQA�s�y��p+����R2ȊTK�Q�:JF�裂V��ق׆�k��@#]��!�4L��VѾ����L�st+�f��W�KB��+��LUn[p�͌Q؈��{r�|���ݓQ�1��U�DH��+)�+&A�(���>f�N^ ���:��3d�f��R@|+y���-;�~}{�"��h���"X�����ח�CFD��\�É���e��Z0v�B�5�y$���=JO!��R�'I5���we�.�I�]6�u���G�9b��ɳ��-����u�ٴ��!�rz���8��Boh�Y���&]Z��fy��U��\�=dQz��K�->W��r����fK<��{��xɰ�b/�YC��y�@嫩���`I:�f޼oԬf9�W����Q>���x�l˸bzW�
�r�E�0�
����3VI�_��^�	���]�?:׏��0��L�6{q�K�2G�B>3C�}`oe&4L���y�@MQ�<;���'��RR��PK��Z&Xv8d^�'O�f�1d�H��y�R*Ƹ4P	۲��E0�g�]MI>�i��R 	5��y>`�g��a�|5y0��.�>Mi�Rz�V8�J�Q���|�.�o��,�����Z[�������{����g�@�L<|��a��>�*qb��w�cJ�8�v�JA����V�#+Wpe�û��Q���V8��ړ��so-@�;��*4gCv��>��*:���(kXr[X}��ex���D�sTM���Zi2�e�Ld��
%Y� ��p�Yq)F�Sv�'-n�ʖ ە�FX�boE	i�� �V�X�0)��	�ا)-?d$��(h`Ǘr���<|���G���5,2 f�y`��2��4�[����	p��od��J���`�:����n�ř)]^���fw_&�+�.��� �s��Z�.��52�Cs:2	�/�F}j�{�#I0c[�a��U��.u��6��8w��PY'B��CN�T7�h:���a���k�B[��LR	�m���r&
�p�9)G�m���fP����u��m����:#�ю�F�׷B� Vx���V���j���!���r'?Ϟ�XX�K�v =l���c�#^q,�:��UƗE�8�	c�?��&t�X���Di��|��^�W6��\���:�qE����!���IA����{���Q"�s�z�	r�T	yP�v·�h�g���g��#�kE�T�xu�VO��y���ȿ&���9LGZۅ9��m��Ί�8ߺ����V��J�B`�V��/��R���̲��=Ы']�8�\����"bU>S���_�I��}�W�;\����Q�����ꬔi�5/�3�S�f�?J���gG���P��<��G@��r��H"ڀ}���R�o"h1-�����S��y-&�i��{6�f�;@�&�	m�V�L��i��X.<��e]��@�P���y��=x�˘�
[ V!���4	;����XlxV64EB    fa00    2bd0&_L84���e� �M�������g���!�in������Ջ��6�PGN������Q>W ���|o��<Y�x�ÿ'��H
�����7�`?((\���tI/���5fd���T0���n'O$�If���7=\�Zjz�e�N)�.p;�g��|akϊ���a=��V���1bQJ�PuX�N.��|��7o�����jca�_�W� �wQ���KY��=/�я��h
��R�4�﵅�Ɯ,W��\C($10?��(�?D ?ד�����>�eUQ>M�  �a�-=������!&�^孭6���o����3����TO���M� +��v/L�Qş��}F��Ў9/�uCbO�F����[/EɆ�ț��F�[���,��Y^~0��Gx��#q5�A� gK'�r�P�����oy  ��.�B��o�#c�ǧ���Q���S��k�0�f�(�8��mB��B�Њ\a&��h�/�����_��(oꂱ!���E����b�-�/�y��D ���ye����@4_��Q~��7�ΐ�����C����U�6RiiEj1E9JB+b�؛�S��q�쁎����MU��;
�,�i_��EFI�6t4���i8Y츱F�(Ú2�ī��쇠�
cM�&+_�)��2�k2�$C�̔Wb�����p1}��b+���8��y���>N4��Y��e�vF>L�0j3��I�N,ʦ�ߟ
�;�6[*
͢J����$N߷��װ%;=js��#	�v)�L_�A�\���̿o�tj�H��cP�;m���F���ƨ�n����4�l���;��0���Pb'�:��W�{H�����N�o��Yt7�	�D� 4�ʷwi�˹�ْ�sE��/�
��jg��%��x(��}L�O]���ڭgXӮY¼�����{z��ap�U���*?�(x^���|���hJ�#瑄^��˷ bSUV;^Xʲ���P����j-f�ܻ����^��ݴQT��|��� a�G۶}O`r�]c(�Zu$��S�f����D�3}�ҟU�ֲ�Aã뙤a����7����2�=h��u��-��zP+�4Ca����i\�4z_6��Bg�M�q�����T��,C��Ri!w��+P#c����;�m�
L� Qrwă��q<��i����}i�1�|4B�4 �(e����#�A D�M���&�F�x����֬�n�b_Z[O�h�J3e�y�h�]�7�{��l�Xi���"Y�j�G6�#�A��x�}�3�ϼ �#���"�!W���Yѧ@Q��	��9�N��H�䷤�����S����$3��'s�*,�b6��,�A}��n��A�#�0��G᤽~�����\ﶔ=�e��8��gV[��I����!�m,6W�Ɖ++�8���ǁ͖��ؒ-M�ui�q@!J|˼����U�Z�+ʍ�=�����zlF�P�Y���� T�0�v27^A��F�}�i��JYE{m����m�~�${J�Is%����88C�H\6��I�X�,��(���p���SI���*�+��u���H �~�坤D|�ç;�2(������L�/�	\�֛�|�"���lΜXAr�sAy���7����)����gW�T��N%n�Yw���ݜ߹���օ�[T�-�iּsQu�\3�>�KS�h�t�i1����lO���*oc�tT�W;��uܜTI�
pY�񿧥�d_љssQ�a0���GTs���v�:����;�I���09��m����n[4p�efs���8ݤ#�~m���TC��r����_�� ����=η/�֓��-�l: �}䆳Q���?Z8h�n[G��"=�A����{cH���뱻�`TB����#����j6����x��礳�>�(Iv��@���Zs|m'�c�$(�n��+�@�`�h;ie�������Mt��i��҇4$��K��:���������u�Ѝ�@��b]_cL$i]�Ͽ�T�p�i�����\|�̺g�+Wf����x��+=r�	�˻�#h�An�W�WA�>S)�ߣ��҇"8���0O!����<�)���gG��G��98�q��P�*�N��{֫,���s�	�5�6AL��^���=mR��5'�_��sE�p��Iћ��7�>�<�΍-L�s[��8���T]�fĨ�K)��$$?x���6B�~�T+U��5�^�tTE�%����~��l<�.Kq����듏��Q�j�[�O���
ghLC��Ԓ|ď��e�51Kי!/�V� D�3>Ձ)�Z2#��N�o�'�Yr�qP��� �!c�7Vb���a�������@G$�C38��H'Z�7|x�;� c�S�~�j�s����MAl��-�gJ!����^!���() v5;�?1�48�0����w$�p������4����HFR �73��hOv�?ˀF3�;���B����	�w47�<t���a�Z�_ �y篟�y'-�QP�8S��s�䝇�I��RkƜ7R3\�s����hC�4_�#
���!��QIYs�w�y$������0�O��3�[��2l�/�p��#�U�f�a�����ѕ�1$�%�>Rc�ǫ��Aڣ����̙���������=��FrW
�Vm(r�!���t��wI��CW`�?�W��b�a���QF�4��`|�����SU��;��[���r	L'��@��u.y4-��;�RC������S�C6��;W��`��-��v���t�����i&�*_а���v,Y�,@WO[��r&�;���3up��!cS�M�BZ�U��S_�k�%�h�eN>@�[K�^]Y����v�{��.}��f��y.^X�^�M���0y�����@�O��-�6�A��L
y�,N�!�`�ȥ���U�9Miދxϸ`�ʲ�2�b?	Jг�P��H))�^'Qp��m��2��@S^b�Ƚq��+Y�zI�~��&j�5:����3�*�d�?�����c��ƪ6ȡۥsm�{r��k����	�r6�Nǆ���^�
ĥʢi�M��o��Z�eJX_]䴠�����н�A�%�`������1��E�z����HA�]�<�n�ꗃ��ʣ4|zxv(�[�|��I��Uӳr�) ���I4s7]��#�!��׊$2�^b^~�o$��n@xn��D�X�N�-����xB�@I�y\G��}hoxieI��ɲ��["���F)0�G�w��# ��oQCڲ]n���,����@E���nf�lN{&	��[�i�Һ��µ�� ���2�{|�S�Ÿe`�����q�q�L!eX�gWm�O��;�R�B�`S>R��x���ɕÈ�b9�x��[�奯�X�����~�5�-�P��2�<*Ek���M&��.9�
<F:!~��L<pJ�ڮ.;�:��
A�NG�b������fl� a
�G�. <��Q�.�H���v��(%�`��;7�G~�/7dT�I:qdNHoC�F��/�^�UT�/�^vǢ:P�򴍆Я�%�Mn����\��y6>���5�Ǵ�c��"����P%4Ty-̽�%��˝Yh9F�J��셨r w�b��1�J�A���J��}�����]�og(�#��L�.<+��{�|�[�Up[]^E~~h͕�m���~߻r�2��p�,͐�.�w9T�8+��WZk��)�_}����@Ǥ;{�vN��	y��i�)������s��-QξՍ��/q��5��h�§�~"
�+��߯�ó/���mF�zE����!�U��<�dEB�1Opt��l���Dw� x.{zk^���9D*p� ���Isx;9�e�
<'� �� YV��=$&����>\.5��**�|L���Y���ok@e�K-z�̯/\����y��s�H�\���i�3��T���ۡ�ԇld���O!֏o*@�졙�?�L-2G��^���
Ɩ�K��\o,ɭ8�K���w%J�
����R¥r��Q�&��k�i���,�ђ�<��M�R�f��'������g�ԯ�tI�����<���Z>�	�5>N\�ݻ�Y%�6y�<B�+Z^�tπ�����U�B��FCE��'\]��� � �!��C��r�$JWdo�"�\j!0^���S���Yq|[!��Up���R�9����&_a�c��T��S���%�	ʔ��; �ɜom��T�`]07�*w_I��u�N��CG0`���1��C3�Զ��%��0��';'-g�L�bFN��  ���YĐ��X��.p3(&�Tev;'t�)wp�S;À<���<������on�X��;^�D�q��9I��"��<�}�\6,��
�b�\/F�ȯ�$�S�ps��5Y.�=j�����ef����F���ư��"��^�E�Һ�ɖV�I�)�Cs]�	��]�]��!�B+c/��< ��TI�RG�W�闹�/T/˞0�v�q�<'��r�7�3�[>sͣ�ʜ�)�Cg��Bɵ�������J�B��S��$�c�{Q}0"�2[�y�XOD�i&O��m�\�TKh���#�'�r�4x�V3	����
sJV��ih� �~�=��Uy(�38oT��V/�i[�ݖU���mQQ�#�~���F�+V�|n�#�����_��ӟ���r������s��5��O ����ge���\�:��z������%~�V!�WBi�ƙ��Pb�>�6̫�-�r�2�L�Hn���<��U����#cp�L�kהּ_�I�>�i�t�$������,�%6�P�n���<�HH25@,lY%��qf&��c1�%�~O�}7u*I�f����dAǁ O�g<���?#��R5?^��L�"��Y�����<��(��wE��4}�10�iIhY�DV
"Y������3�%܂a�ko��Y�Eɜ�|�tnh��g��'����A)��.�*��t�h��Z� �XHޝ6�Hk��c���yy�ˁ�$ޟm��C��$Z�?���*o7�� ����X�d�J�8'�R��j�?�U���"���o�����*	��e�bp����6h@UKy��m�j~����U� 2��f��?���%c�op��'f_Ԃ�n06$;K��a�x�7bc$ ��ރdJ++5Y��R:
�)L�_�<NB4���] �p-���C�.'��'�"~P�M�R�b�˳ӘC�+�0SAKx���'����Ŕ��1�$|0ds�Xa�E$q1H�.ej�UOo�&o�0E�tX��kإ �ڑ�����vmQ��;���;�F�gЯ��%B?�Qr���.����z��+�Vm%�q]0���LN%����
*����1)[��>(w�Hb�t���knى��ä8=2�����H���@�,��A2����a-npY�gkvZ~,�8JL��B�m���� ����"tr^�+���&�!�`v��U��SфvdeiL�M�8|���g�Q�?��υ)~�-�?�^����"�A��=��	�Υ"�ʛ����V~���]g[�/q�A~/h�*��+�i�7:U�I`�a�+m�u���P�Տ�G��5oQ~�&)l�l�ź ������T�+���[)0N!��a����<׈P��۲�tZ�8��k��yO�R�l�Hq�i�db�t}s��l:Z�69=NfAR��)Y�~r9��*Ũ	�rs�s����#e�ϸan����4��NG���qXQ.��'O'毀3�i3�TEd��Si��o����Y4ϠG����GE[	�	фh���	��� ~�%�IF7P�Ô�.��oǎ����M�[��5�qƃ�rځ���K���W2a��C�����0�]�,		�3�AL�+�Ǖ��[{Y��4n�g6�X�碀 ��Jۊ�Pf�����\�h�߲J5�o谙܃m/ �Pͫi70���``&�s�g�׼y*�����!�C���HT+9}F��iI�W7��[-b�^��W<M��%`P��$V���s�t��^�Q(V
��%�AM�/TJ�
3����D� vސ�D��pi@P�2�1�5�0{\��>Ͼ\�q���b��^{��cl1G��G�q�{���q9s,Bt���k��Q+(#�x5:Zծc˧b2.�kQZ�	�!N�i�n�7Ty�u�I�]!�\��ҧ ��*z��ಬ��GS8\�a����KU��l�/rd��2D��i�x��?�fS�}N�+��s-ǋ��P(�k��c�Ოoc�6 fNQz��nK�c?�')��ܤDB���d�x8o�	�2ਮ�U3*xc)�-���q��׉R�����c��׾䉳�m��SO�ގ\�>+�	�,	X�g�X��a�X¯ׇz4�`�uP@�_�G���'F�S��lm�f+&�}�lI��H���f����(���ӻ�u��i�ֲ>N��y��� ���°dO�������s%���d�/����rA��phN����;�����G�Ba�nSL�j �߼��<X�h�P��!�?%$M�qu�\�MÔ�nhd�1�l��#O����B>А��
k8;W�+�9��r�k�<6yFAD��eNNEjvE�)�Qx84�@�Ԏ>�G�����g�!h���)�v�&c��.b]����!^�q����Fek��y>L%-`h��z�X��Kg �DmVsa�G!FBܓ��H�2s�q:)��U�Z�{ְ�>�ȫ;�����$���?�&���0}{�j���ބE89��qh�"�{VYX�B��I��{M�����d�3��}���r��ҍ�˿q�yz�q^�.z�9����y�h�S�w�Z'}�n!��V��T�c�`N��mv��w����Tʸ������qᅷ�8;v�ͅ	�&O����.N
�J����$�(�(&���ɕ���3�BjcH`i��g�X���ZQ�D}�+@%�R��.�,��Bш��c��T g[�4��d�m�|�p�i��[�߃/�wQ9^^~S"^>_?u�
������u�$k���N�~1�p��i����f��ɐ{�r�$񊨵�l��Ф�W��V2��`?`G��fu`,���-erօ`����j�&�UT����3_�ϯ��҆Y��ig�r�i�@$b�'�؉��KgM�g8�t��'���Y���hns��*�\�\.D��V(1I�F�ۊ ���7������DqY�K��q}��N��ǃ	���wnAR�D`R���/fyܑ�ȟ����}x���G?���T{!:5H���TU2���������� :2�����j�u%�׮��-Q
t�I����}�bܬE��ބ�����Z@&%`6�&��^5�	�j\4H�qe�=#7:2��/�d���9a}<pS�Ȝ�)4B�~����M���L�?c�8���Ί��pBP&RE*��v�.�ΩM�Y�"�b{��^?S4ԬW{	1UҁV�U������Jj�nm� Z�h���:?M�nO2q�:ktcf�{�$�zm�pm���Q��Sʄ괃���荡,%C�쭁Ȧ���0pG�v0QЫf��Zw[OIR�Q�˚�/O���� ���_����2�A��X�ZT��q��� �=U�Ž�x�͑]7�v~e4JL��eNYlx7Cl����V��97����--�~�I�^9��f"�,\������r�ݗ��}���R�oe�"��)�+�����AT�䃄by��.�%2�"��k���߽�Sbb�*�H3����ų����	����4��Йb�i�/����?���y�[�J������Y��5̷��nҞ�g�&�f�}��<T�J�LJ��sz���FPd����Bً -Հ�sl�j�A��Mn�z\69��<�ܒ!�Q�s���9 � {v�"|��`�CO�F���~n�m(���a6��l$H4�
���6��T���������$ö2X쏩{g������'�]�t����1X�cܤ`�H)s���l��2�X}�a�;��2���w�L��,�W��! ڵ�v�����5�,�U�r*�����ڙ�O]e�N����}ƅ���p��'�˜��{���%�C��Lw��M���ρa$��ő7�in�U��L3?�сqNd�g�'&1g�]�j�zP���Rd�ua7&�!U?�\t�aJ:,��d�С�5��M?��c�ȄH�k'�Z[LZL�Y�`~�f�!d���t.�]}���͔��M��.�_\Q���S.�C!���H��e���� K��b��k���SU{bQ����!�V��-V�?��Eu��zS�caҍ��#.�Hn� 
�>�+�	O����?����@먁�/E�>%ic��X�0�Ws�#�-G�]������8�D�Ѻ"|f��7"S���Z��|�Mz����6U6ql� �?�x��Q�]H�G�S��F4n�fy���*���آ��r2���ݝ�}nv�XG�N��L&�OY��~�?�H,�uF
;�i��sӸ���3r,�`�]^���;�ɯ�Q���Ђ��e%(	�jS�Lk��2x�UPع�ؗ�!؂�������� ��ꓖ.��5����>�ud��'
i�����m{�)G�~�߻'�!������|��y(mk� c����Н���z������)AQa�3�C�Z{�����8xDW�#�{j���еd�|"�ysS��`�xŨe�F1��,�_β���O�1��>�J��:\���da���������1���E�"
'N	|wqB�ȣ��C�׬���g��r ?)��Y�T'��3�&ܧLh&��\ݮ��Fk�E�c��0��0'.Ƣ/#��F���݇{�eKwC��Y�>qI�	B)K�X�PhE�����J�Y��y�B�d7�).Pr�p%u(��a��B0�[�5��fcQA�!�c����?�Љ����n����'�Y��6o�"�#�93�N4}ˎ?l�C��J=�%e���9h\������1E���(�2sz�t!R�b%p|�Y�1�pHr=�$��쑟ӆ�j�2d�X+gr0h�T���N�Qs� �n�h�,��e���r�a=��7�Dq� w�qJ`M}u�DRY۾�]�֋|iv�r+�*�0��m�5��_,�9�H�!|�u�L��iQ�!����Ʉ�b)
�Z��1��f�ݸ"e�[��k�>���G?8u�٩�(#�1����7b������jZ��-�/�*_(4[#h8�.��)�#;q�=7�mg�+���� �&��NM���(�
M��u�g�_��yQ��&��
��I]�ح;�%���ݿ�/&Uku ��*50��qJ�=W�V0��[bT��"��Ar��E����8�3{�nd�L�-V�&�?������-�-���L"�K`�T�\��-�>m GSH:���w	�Z�I_�b�'�=�L!�U���x��Y�g^�7*T��b1q��b��/��I�[�$,����9�SթȰ����1��.h��Yf��"3~����m�����i-�<ŀ[�v�FK`��%_}��/+g����cr�?�|�[�b	����t�J��ށ��i)!������#}�{'�)5u���X^�9�24I�u�$�*�*t��	���=�MѠ�0x~��� 7��&~�~�����{}������ķڧ!���R�{�Sz(i��ڋC%�6�`�up���E���
 ��vRq��-�_�����/e�|�W���$��.�r���(/rc��]}>�6�C�*�Y�PFCmO�ob�ɂ�R`M��/���eNpC�G7�_q�!�$Z��f3e������P�궁=��4Y�A֧�w��qώ��)�v��1��'�l��������x�C`�3T�%�>�R�+r�zH��u��a\y���> �:?]P�(���yC��]�1T�Q/��WL���i�C�A����'X/��,UR���̌�>;P���#�_�]\�$f`"�LA��;x�u�x���P��nhl� V��e:p�m�b��9.g ���H���(� �0��h>`jx	�Z'�UN�i�, F�j�H��
β2fu�$�сc�u�����b{��D����Y+��������M��|<������
���-�/�Es���2F_e�O�U����z:>�i���CU>�����E�����x�J@���J5�.o�e�����okX�q
��y�L���&�Um)'��%�A��\i�d)g��V�?.�ٿ"y�i~��^lq?av�e���n\ρ��S��Rl��D��.g��T��f.��dl�5\�.�����K�.4��hh��R�[����c�{1m	9B>�Ӫ��6a?���^JY��	3��[r-wx� �D�{�ݩ15�#s	���M����4�e��|�������j&r�"��<%��i���x]L����.��3�P��M��0%1��K�����Ϊ�v��س�
[k�!�-�	�/�לoE: �����i�i�fq�)�]�V�;�x�niA��c6Բm�N�C �M��ˣ��d��+���Hz&5�7u�T�@ʤ�f�+�����fùb*�z������4�]�'���*z����m��Y�
Գ�pF���HK	�Fm���naw���V���(>|��K%P�&�������n�G?*���Ny��l�_S�h�.�N��ͺ�q	AƱ�
��,'?p?�ſ��/�ܦ܄7B�D.v��zwZ�\��<����x��׿�B싧��t���vU��ka-�&���,��5��ǆ�6A�'m�E�V��D8gT�X�)-�+�x�^�}�rn�o����%�Tt��p���DO�Ә`�U���IL����Vp�i�3�w!���i\��6�.%o5�$��k�mWH��NG�r��(m<�:�f&_L)�V+0T�7�	Y���jc�5h������e-M�Z�����X�\]�>S�Fm�ߩ$�w���^���dZ �:��fu�9#������/L)È4Q� ԉ���ly�}���XlxV64EB    fa00    29b0��{Ua�2�V���;�DNt#���ˠ�����Y&�$I��(8�5^A���+ګ7�R�n����ZR���	?u�(��JA%�D�츒�T=�ƶ�n�Ô�[�y�,+tHv�BGε.�@��"%��F<�l����z��}��g�x�:0,>cK]/ �	�khr��A�xX��HK�I�^2��^P7��<n�*�M�����/e���1�X0\�<��Y��K���5^�d?��Lܼ�%4�q�G��Gx�����;w�2�-p>y�`�u��9v��nyhb?*�~�wW �]�p���P�l��o��1_�,�w��,w�3��|�v��sBy�q]#��o|�C�i�~���{Ӷ2�_뤫z��G5+X�b5�;��[��i�򟤡g%�,���- ��ힽ�y��_��#Y@����q�_�sa��N J��xAL����Z=�����x�<5�S���5�L��V("�v)���I����������Y�^�X.}����/q��	E]�|�6�!YF�@��?{}?J��ް��$_��p������]���|��{�o�}Q���/�����	�_�K���w����H����+���!𢆪s>x��]��i�a%�9Q�wGm2�-��I*r�ϋ��v���*�Q䨆�
�2k��&`I�?ˆ�Ї���� �f�PDX2�o�0H0<	��Q}�Z����Qj���6��Ɠ��x�ϙRX,�,���[�&����,�P������_v�_�J]2=���vGpC���Y��.0�*��Q)�4���n�}�{m:7����%Ď�d��_���00�d}N����H"�Q�v\S�~$�ѣ�`�����ʗ>"��[�b�\^�t�hIN�N4<����M{;}k� �aQI]��ވ]A»�;�E�0�of���mp�f�J�)j��D8w��j�ԍ�$�m�{������~�7���>���=��[��33��[	����]�l2���}rU|����2]$h�-� ��h�����[�o~�>���X����m�!��0�����v&xa!Z�\��v>*�|U�67(�x_rs��0�O�����ݜ�/�q�=_�RhK�&���߾؀�Tݳ��3��*�`��i&�/�U��֝^MPI�g,7�B�j58P������JYF8�+�J���)����Z�vw��˃gW��ܾ�t�����"�^(̸�.�Da�J�2��cE��>���Z�(�iK��UM��Gy"�y��§ߧ7���{�tU�}lo'�j�
:{���ͫ�[��q�%�C�AuN��1���M�܋���郤g'�1$F���������2{�т�Ңg\�tԇ�O���uY�3^B�WM6��_A�c��W��Ąt���Y~�z�0���hBD�K̜EE%>�?K�uR����$���f9�o�+$�����?�B�T�_����\�~�1-�͎z���X��jn���6xU�2PM3��2n-��k����3	����� ��ʍO'��׎9L+��"/����pm�U��4�K7�}��^�:m=�Xc/���M��דr��FP�|�( )��Q�W���T6��'j�;)lHԕ���mm�9Xb��J[�N���D���o[}�@�f�DG�;�Ⱦr�[�8u�WU{����7J$q�ƨv��3 wc*=+����CO���r��^m���ڍi�R���ъtΆ��~�>�#�8����[A�g��Ս���F�M䡥�9G�N��.o�XN�ѩ^��H�n8����cq2���qk���>Z�^��_��>{�`���)�2�Ɛ�T1�
O�@Z�s��c��������j�r�7_C�~���"Te
j*[�*g;��<T����򂅦�5g���VV�G�;)E����S_���X3���ϛ^��-!U�$ߦ�HJ���v�A��ߨ.�2���B+U�r{�J�Q󅲱j��k��\jSU����<�*2�DQ����D.�!(d0*Rg3�	dp��E�|�M��IN��J-��a%�%m����|'��������G�OY�9��iK��T*k���y��@��v��q �%\g�k�ў/	Q0=[u���~�Y;x}����e�39ǎ��V�:�E&���H�A[��u�2�R�y[YYg&\P�J���e�����ˬ4V���'�f�̲��"؇.�l�P���n���t�O��Bۀ�`��m ��>F�VJ�j��J+�1uu�#;���v*�Y�2-}���C�m�Ӣ*��hH�3�1��r:�y��L��֔1�Z�1�>��Z�S�h��RO�CxlX�5M��1�é�>��ڞ��z�m�.0)~�(�&.�O�z���B���?y�fH�9s�z^����-!��=tV�����7�H����o�_ԇp9��~��߁G���W=��oq ݖ����U0s���T#$��Ӣ���vM����v1�����}DAX�����6�6:A�l}���
�:�N*�S�_��vL����c�ӭ��X���Q��A
{{^�djӧ/ٜH�8]I��+佤|$v0e�Z,�^➋������:���}O��x)W*�}	�K����`/c��d���b�_���B;�j�wү�ҋ\�k˵��k��_��ue�U R���N��D��{��I������.
�[�~������Va���N���+\�'( C����l%Z$����I�7>y^+y�f������|ε��I�X�����T,�%9K�d&��]ko�LĵVeօ���k��v*��c�|=�J����S�͎��e��)+�>��� x�<�����%]T�/7����qTN���5lT�]r�u��=�{_9 ���z���G�C�4RB���mn��r��Vڻ��}g�����S�Pc�O�]@���������|��z,�����d$]��}�^^�����c4W�L��k��7v���q���n�`>��窲mE��H/�=��X9�x�O��)��)9��9� dJ��&i���(ǽ�g�J��m2#�q�|�Z�y�a~G1�0s3wޜ�P�|tb�H��$�2�͵�U��Vb��Ԛ�햴-���ڬh5YP�E�{�DAf�s#E���2�}:A%��x�'�	���醌��T>�~�F�Q��\�L}]�J��^�&z*Ǿ&z��E�VRM�����x�I�S��� ��KOrLP�8���W�Ķ 4�C4��%b���Q�;��7~.�x�#W�1k�DG��v߈���MW��d�m�'V"���$e�$�b��7șB�E�P�o_r��	N�\�@��]�yЍ��Z���5���篸�� oչÄ>�3�6�_ˉ�LS�x�� 4k�_|�{�C�Yd:�1���z����� ����1��Z��+�%�"�����a��s;44�*:p{nˌ�6+D ��&�0����*�F��]�
�e��ڈVmS���pQ�עl�m�G���������K����nʳ<�E��p�;�=my��)��ޜ��E�A�<���Ե=7��Jj�D��\��濡��}
nLe���� ���n����i�ӛ���J�e���9H��+�A�q��Ҏ�z��z�9�.;0)�z��~�pX��+����]�۪�fN��}پs)�T#7П�%Uju�GȺ�ٻ���͔IR� 9N
UDDG�E��q$�f-1sG+�st��,"�o��$Q��kl=��F�^��+��$��P���d�2��Σ�`��퀔\f���>�Ӓ�(�)*��n�ͥ�1�C�*Y&f{��CV�E�Ԉz��,h�_H�&��Q���g���}I�az�K���۝ՙ��;Y��̛�:t���s�Q_�(n��ΌW���v����)�T�+-��c*�z=�!tR��8����"��A��i���8����&E�I�E���r?/Z�-lZ�	LgD��73�<��d}�r  �W#W9D�B4����}������~�������N�y��ܩ�:��E�l����>9O�d�D?�h�b�ɇ�c��<��k;*4$�u*��v�c�����s�*���+�O�����V��"�O�0^!�i����7����:�S�"�1N�|�� r���C=W̩�+�}�#d��⬤|IUp��MN�C
�!�"�{�J齝m�ꐳ�/} ����ƨ/̩4��,/��zӪîe���ҵn��Ų�V�Ϻ2Ȏq8)�p��/D�YX�Z䶆�!�����-���Sc���pK፷��IL��'��G����k�\oJ@��YVrwHߒȍ��&��*ې��P��i/�a��Q��a�	�#oզ�������ʡ���n=Ip/17T֓�9LYPQ��ܡ'C�#	X�?⿏Q��Jg��L��|U�����ݖ��h��}���I�-C��+��Hj�$#��)4�?8�? g���f��V� ��0�I�|��W�0n�2�*T�
�8\��a4
�2G���?�"�Ts�cd|�F��~�{�]y0֤�� 8,'9����s����Г	9���ϮV}IE��sF�)�賙�	Pv�I:t2��;�s8IS�-5�j9����e�n���n�g>����ZGc���� �bOZ��׊�������6�bM?d�FPc]�"�yx��Ϗ_�7�tg�ʕj�rq�L�_�0yƴ.ED���}��|r��Ô6
[Q��8��g�k���0���r-�:���GT�I/XY]��Qr��)�ݿvY�w:4ē�zG	��^�ؚ�f�s��o~V�ք�<�f���y��%�XJ��4�W����oʷG1�JE�7� �5�f*�R��7R��W�"�H���q߃v��,�mlG|��1�{�vً�&�U^����5)?ˣm�������TW;�����;g�K�]��G���7�H����w�P���\�TB�@����Ѣ�L� ��6Mc��o�8N5ubi۟_m�:���:��8��:�}�E����z)��Q6�V���T�����ֱ[�󓼷��F�0��)��c3v ��=��1�%XK� _�j+W�pl��񹐚Ȝi�\ڕD�@G�ǧ{f;1�L�y��8Y!���G��5�d\�y!�-�O�FU �%Ro����J.��0蔰O���� ���"�g�H��:˦1�#��^}�l�4���^�����Ak��o���#���âpx�$�S(�#b1���z�|0}A$����7((5sC�v�y�̶����UϠD����g�V|f�����Og�1��hӀa����( �i��)�T������<o/���[��X�􈵨�㍒�	hwr�`$]�v{R���}a���F3����>�k�w[#<�c��(��v��6���<�p 4�}���z��q,;��짤�]�T��tÔu��J0E#��p�e�bԯ��/OJ�i���j�����z��z2.�Дf����.��\-��ko3&�+���u��Xw * ������M2,/Aiu�Zؘr�uQGj�����˶Q;���M�9�L�&b�Ttg~`�	VK" Y�2`���|6P7C�5��G�ڬ-�h]�q;u�9�6ޭ=�p չ��{s:�\��޴ڰ�!��uN�]�,��u�fe�����H�����*�Z�7]��N�� ��Xo�ޠV��p%7���O2��<K0�|.�kf6�su�ұp¡f�	��Q��8�	]?����d}�U;G~�:p�A�$u��a
b�3���K�5H�}~�2AB����60�% ���}+���\	Cx���qBNQ�;�7�o�����n(�t�䕋 I	�29�G����/����35��S6F�MN��Ums��Tz��
T�mm�_�2W�.����m�0g	l�ʫH�����_s���,���`�f�66�L���{X7�e��Ǹ�"1�/կ�Z� �WF`�uWyȗ�^��H#q��Ǔ���GH1���[xp�����V�yۤ��2����`�
��i$������w *�V4:��l�T�j��AՇP���;/Ag��j�U�|<ä�)�_��g�s3ىh���ψ���>�����Rߒ{�x%�Qq� ���vC�{��b�y!&Kf�Vɝ�Yck^�%#�<�~y��Ò6K�P�z�W��/ ��m���f�������|������O�ڰ�S��!�Z�N�\��{ן!������"4�E�~���F��R��x����e.�Ӂ��y���m�eȇ�lk�t�C<a����SB��V6�>H�T˵�_����)-7u}�Ƌ^��.�޿�LEä@6+�!<֊�^@q���ն�WclIy��=��#��F*�/z���T{��%!�������[m���ֺz�]�5�m2']����QU��3>s�M��C�⸑�^l�9S�?wF��E�#k"���5o����~��܇�#�m�D]ĕ_�����\��4����)$V���ʃ��Q�+;o�L�5�?S�P����LV��kp޹L]�l���5Z�"��:x��E<A��P�%��ػ2���4r�*���+�w���[��c!�6��n�HX"d�O�������w{3�� I���ɋl:���Er�_)����p�c���:N�6Q��]Uĸ�@=�Is�z�뺝�|��5�&M�C���iy]�%>�p"�;�`ֹa�!ZP2,l(D�ުc���$r�xX6�-���&~k�d, Ϙ@�
��$*�0�p�r�%�8��l[���~���F���7��ܷV�s~����6��}�K��m3�Ê�n-v�g�VC<+#�^}�G�zuؽ�1vL���<��O�j^V	m@�����P���q6oJ�]]|o�����w>%�3��*|�;����2_E>����ԃ�I�!���"�����J�PX�	!/2�*9L�\���,GG7^�0�b�hf_�C��xD
�׹�J��07�1�B����*46�$� �X�6g�Voϑ�XV]�ZR9Q��t���8�>G-4�N���j 6{d�����y�Q�W�U�����A�v1t��V�6���`;�*�5#;,oPwX�/D�	o^@����Z�Fb
�^+��B	h"a�Χ�\8O�g�H���@(���q�đ̤uO�i7�ԩ���/�jEf/1[~�rL�n9�q�+�W�,�
��n9M�ތG� ���=�H��*��c�[��/܅�*����F�0�B��{ůF����Y�v�o��F��PS�򬧜,s
��-�g�6���B���Ӑ�۾��۱OYE�R�I�.��xG�:;�7�#O�U��S!����/291)EEǆ��!�90�e_�׾I#�6
�/�^��r�]H[�(i΂yI��t�	��j�#H+j�ۄB�h��7�j��Eh�Ш��g���q�<��T�᧏���z����\���O�_9h<U��dх+�u�(��{)n �ai��*�wly�ǉ^�I����c��w5qsk�z��V��KК{ o�V�3D��)�'�UK��h��ib�����J�TA��p�N���/Sw�eOq��aj.)uC}#z�d{�'�Y�lN@�	F�����<
/Q�g��Yc���8ZE�N��vC���������A��Nz8bVkpvjE����4�7�?r���n�cj�B���A7�V�k�xG��n�!��z��Psnt+b�4Ƒ�1�����De�GW���C��SӉ��
t;NF%q�B��}P��aN��$#���/�m�fi��X2-'�떎��k2#���k��\>Y:���N�F���s�Al����:�G�(���� �� �
p��D��+�8��lp�#�jaȟ������T�O	8�94,{#����~_@����½��̷��8f�{kb���z����G�5^��R�.�(�
��@$�;�����]���P�A?9�s��O�����.;��S[�G���Ba��ǿ����[:��9DP����JT6��#4n���˓�J��K�S��DLi�(��^ൊ�n<�����&.b��2PB�^�I+�G���8z1#��Z!zB�>"qu�3��DM<�љkm*�C�#Izd8E�#%�u��ǲMh�y+� �0 �ÿZt�EM\cN�2��L���Ue��mg�l7����$7+�=7>�{�I�g�K ���.�0E`�7z^#����3K����[>7Ii��Yj�BH��Q�,��WۅD�D�*~y\��@�I�؟8i=�NB�k(Kx��(a���2�L���%���HVi����^qA�*)o�X��i���m#f͘��*���5�Ta��Z� �&�b G��q9�4k���?�TvǝdE��`tm�����H{ �X����e�Bs��ɫ~<]� �}��\ǽ�Bl� �%c��1��l}�3�P�=��AB3��)�H�D��� :�|o��u���h��eݺ��^����W��*&}]��1��i+	�_�tF}�ܩEN�9�Z���U���S�=�H�3��6��c�媢'��튺�IeG玩�.b|A. ���m�v��t{p��p�����<���L�Y!i�*س��[�}���H�D��:���y۰�av��f��8ZA���R�cQ~�d��~�&�GԢNp������^Q^$fX���2J���;�U���6-Y���?n	��	�r=����(��u|0F����amV�y�`��W�~���&"�z��ꇉT FS�4��.t[I2,F��7�ζL���X�R��^"d�6Ũk1yJ�����p)B��aS�ge}�H�Rz��悜���;�M[��QR����h\�������W��W]Q�+g�'�>X��r�ЁI㯛q/�h���{-�n�He�q�D��.
_���,!���J��(������+�c��q�ɿF:�%r����FS�M�B~�鯏r[��f�@M���.�ETpo�Ջ[����\�N�ݯ/��/�f�R�Хh��#J�3II�r���)�h ��e�:#�s%�
���=�J��X�Һ�2�#L��#�����4��Q�O�;\��[.C��*J�9�����_(���*��XI;���?��d�Y�<�#�vU��п�@YP�|/.8����ARۯE:�N��b ���x~��F�c<RƔI�!}ߜ���/ǯ��NMN�d��r&	$�A��`�<JWC��R����)���݀+��(I۷/�}����<�QV�>�ɔ?15A='��"5���Z����;�=�lMZ�fPR@C�l�K��L.*h�҂܅�8W8zϑ��xK)�ahK��ۭ�K�2>3ٝ�޶�z&m��?d�ȸV�ra�a��c3�!����p�%^^Ác�ݟ/�N�$�dQ""D�w�'sb�<w:E0�+��q�d槟IY�����E�]���G?z�M1q��1>���c�1��%�w��*&�o��m�C������s�\�Q4Rɣ���@�&�
Ԁf��?�ȏ�r��w7/&�t&�{B��߸/(Y���������H#��쒭Y��a�;\��-	�P�Rl~8�
.���S�8��B~�l��E��ݬ�6+>�Z�K%�Ӂ�n�ғ^YQr�3��6�6D��1/O�( k�Uʸ�]T�Ӝ��69�ؤP�\����Q/��p���2�v�9���C�G�(��8���1C�s1��"��\��� ���J@�n�2��0f,7��$9�њ��L���J���}�#���f�����s[;L�v���ئ��o�׾�r��������7�����ƣ[��p�~H�d~�k���LW�ɡ��E�"�5�E�+�|U����xD�Fܶ�UaH�΍g�1���Z&9N%s�&[C.���˪P"���>���ԍ��9�u��;��|b��Dʬ��9Q�@����!倓����>��ܸͤ>��(G?�RЖ�x�h�(��',-y
"��-a��l�Ƌ����U|�<%0Jdm�$�^�!/�^�	��tC��Z���{WS��cF�`���T�ZD)>B�ֽm�ZЊi��Ĩb8��ߌ�t��s��5��40w��/�d3wV�l[|��D��ͳ�|�a��.���cF�y�����&�q��ZH;�A��2�+��J�Z/�VrM�<��	)��[�|��ͮ��I�QT��ۺ�J������N���$�Ǫ��7����|��0�r�+��)HmnF��gB���7���#N 7�o!��É&�qn��{%���F\:اU��F�!���J�b��#<�(�ޮ
�E�eۨL����)7�s�Bm#� �3wI�@�U��VY�+_��
L� 䲻&�Bl!oCM������'q��5��$�ט������1�}��P��ۿ�"�:`,eiy5��V����X �a:���F�'���7^$Y�3(�O��^��ϵ-*<�R�[Za���d��?ݫ*=���H�q-���Ž��ʅ[-���XlxV64EB    3424     9c0�ߥ���ѿ�)��%�U��=N��M�LK#���4��yKcW�D.T�.�;��� ��o���!�<�~�5U�uԺ)�N���.��!�l'.�7�d�� ?p;P�:�6��pj��g�����6"���$�x���Z�j�xR�X�w�Q�|�����D�+�U���b�v�T&�xwCSsi�ی��;�y3��Ce��|6nsͼƘT�*�	:�}~~AN��_ã�ʊ@��eu|���@(�5;m����U�b�v�L?� 91�}�`�Q�#�\����;���:Vh��{ZQx=�>��nfC^Hok"?��o��SY-=ɡ�"��h<?�"��o��=c�7������Qy*�ԃ��N�����],E46����@�4���Dt}q��}��7/�Q���>�(���e�x����_��Ϗ����˅6;ly1Mq[8b���Z�(>��~�9v�����oC��m��K�?�cΘΓ� ����y	�kSb6u��u�2���A�������3ݾ:��|#�c��Ǳ4�>w{����*�U���^ �u���w'�^YH@@ �/�'�T)�1����O='Y>ZFX������S�@�M���%�.�<M����ȑ��Y�j��ITdFc���<���k��`K/D a@J��@
��1x��q�P-�%B�GF��� y?GMu��`��r�@�hF��V3�Խ���13r�4"�TQ<�B�t��l�x�Fm�7O�I�mm��<e�ɢQ�68C.SH��y�~��`���5 �|�0��t'$�g�""�=���J�2�0�٫u�/��ă�#���wCD�I0T�enn���g��1)>��U��b��@�9��Q2p@���h޻�.&?�q�Z.P����Nҟ����>D̓(���a�V���+..�V(���B&����F�a#�:Ș+"�h���Q�*,B����D�Kmo�����S#��W3q��_+J�i�]��� u���h~��\}y��Y|]���7�n76�w R� �Pς��r�j�ה|�I��*T�,Mw=Ir�Q�������2G�Z��<�x鉷��;g��
��Q��W��[�r6\}Lݐc���yF�1f���#k��o.倡��`%rU��0���5�)�e����#���Y8͢P`p���Na�?��� 1�x�@nIM�����_�7f>H>��L�s(O��G���U��&i��&'��Yև�	Y\��Y�(m�{=ѝ�J�Uݥ'�b8HUP���V���$��9J�(x����z
 ҋ��Z���z'5}��__�Wrȧ�S���(C	ದ,�������g�8�N�A�bW �"f����a�BL%oo8N�{��&0ö���>-Iȅv�"�$/%u����\fIK�ʱÑHL,=m�/�`$�Z��5'J�jW#����(� ����$ΐ<�b��9�<��F�/Mjֹt=�Ÿ�A��UʎQ�%JX���Y�ZU��6ɠ5/u!���6ۛ˘Yb'h(�{t�����ϑ��뼶M�I3���b�V��}f=�3�KJ̾L���Î'�d�C�Il{��v�{�b���)�!e���z�V)5����Ji�x�>wǳQ�ٱ)�:�,7���f�iV+�pZ�1���H��/z�Y����,\>��Խ�@���>{���<�(^f���~��@2��x�V��.+v�߻*|�� ͢���Ee�J ��9J�]DO!n�}��ųM`�3AL~;��Ź��<J�ƕʤu�=<�����)Mn��L����BA�3pFV�Lg�¬�3u+�ws�ĥ-A�'*��t�z�ʊ)W~C���)Mey������׳����(�+���8/\��i��2�i�ڹt�a6�eY���K��;4T�h���A�D���F�>�:�TE��^�eD�&���;d{��n�l����޽��Q��챷ق!�6{�*l�(�?Z{?F�]�*��G�j�h��&��\��vi.bu�Y�d��� ��Pqͯy���o�E������:(��Rү^���cS&.Gl���{6x��r�.�9i��ଉ���E�Ʃ�>���$��F�8�DU�7Ŝ����|n93����mBS�G#�7�S�3i��(!�c����㥍�6��2�_dz�"��/*Rs_kィ93p�N��\��4�(#��Ds���6���D�8��ư>�nj��=?Gx�1����k�� ��P���v��{ )��	�?z�2q�	����WD��5K��7���]�P�3� �wK�ڒ^�Ÿ2T~YP{��8q��Л�K�t�ĥ����$4�>is��S�v�ü�9����0��L�[�ۻI���[ڎ������.�0�=���!�:m�$s��1d�[��C>��j��|��*���8/(ށK0?͹��>7���]�q"���l� ����