XlxV64EB    6329    1730�=�ǊF��,��Da�� ����A��'L䭟ئ�Ӂ�5&�-H_���;���/dϿѥ27�b?/;���=�鹊9h��I~W*���J`��J���tR���&=?Hxւ[Q�V�c�8o��.'��(M6���A����z`7(aI�m�^�齠J�!�e,ƀ���dס�ޠ�9<_Mf��y���ʲV>|������*�)��������4݂�gԴ�AN}�`��.z�p�%X����"��-Xl���
E���l��<�F�T�Ckﭙ9�3(���.�q�Ґ;w���[�Z&�L`Ԇ�.�c��'J�s�}�s�W�&X߬Q�ë�V�yYX����h�x����)���5�!�aS�8 � 1'j��GHC���g
w�ҎdT���0{��5�{)����<�(<�/�6�0©d�&�0����P���0� ��t���% �������	�袶[=M���@�Y���Ƶ9��:���v,���ӹ��GM��h�~� �U=Z�����q�ݢ��f[1����I����PF�id��Ş���{q�7���y���F�
�f+�r& zu|�Γ$�P���H���oD	j�E�EY�?���<=������g�#�.�J;&��7����(`JV�-��LS��ǎ�<��=�ΌES�v�w���z��j$�x��5$a�G�Q@Pd[[����Kt�Ms�M]c͒��T`��'KF��)۞�8|��.���a�6C�8�Q������_W��;~>�a��X���fI�6n��˂��Y�7�8pZ�k��z��b�_JoKuN���ɿGjv��'l�:�D�X,'E2�}r����*+c%㢤a=��fTb?	�ÏX�9�Seh����SKF�R�3~o��:'�6�Z����-xJw��a�X�	�a���,у���@pg�yi<��;O��	Ό�P��L������cb|1�.��;�\(q��o1Ե嵁(��q����p�\��*�G1��Y���ot?7��ܚK"�)�1^O�i�#����Ip�c\2e隶���u�Iz�O@���O�ML{��i`� ���~��;�m�t5�U7���,�䏧8"�G<c�XO�l_'w�zS��el�g��X~@r!,���OV�Kr�f�iƃO2�1�Z�RkH,o���K%������/�]c��F��=�P���;��OI�����&X@����"э�<�غ�|�%c����m^����S�1��O�-ذ>�yp��Q���0^���1�&u�Вs� -.|���a3�DDo�P<���n�:�ݘ['W[���W`�[\��oI '�n	��5��5a�dc�� ��#X�!W��^��j��E<���)ڋ�5�K�� D2iӫ��#�6�ϥ��Q��<b��uR} ih��y	Y�&�x)�Ǭ3ժN�!3�}�U�m���^�psP��U���z���!��z�mN�J<.~:��]�y���@#�d�T�:�	ڰ:d� �/-�5~f=�.��̫�d��Y�OS�+,�F���=�٭��
�CT� ~c7|�<R�dJ�[/�l
��k56a���P�Il�����K�2�wb����Off�#4ؑ
j���ϰ9X;�IV�2\��S��wD�@X]��W�m!�b7�̸%��X��-c��nd����JIA5K�M�e��'DW�u{�8�4TZ�U��UV�d�7�?��s�'�}ܺ��p����Lm��9�Ϝ�*/,����r�g[�0%!��R��� 2\�����M7��*���7�p�X�|�Ep��G[��Fmj������2;o���G�s�����)rZ)�*��]��)t�g�=o��j�"���gu�|�Z2�o��Y��'O�e���5�VE���K����>���E���U��:����"�i��M��ÑJ�b%mJ%4�g	�f?[���X�	��\p7��=c�Trl�h�:i�-k�>	o�|��v ����IY�@�fh�8�@ �pa����o����wR������.�?If0��6Q�qJ*pAQ:��9����g�0��˼�(Q�~����j���4w�:��J>q��-J���lGl"�7� _�W� )��:G�`�Q	h�Â�Q��P_����ދ|UbZ�%ՍYi�V	�����f@��6	���W���hE�|Z&h�y*�eUR�^�/ �pI���>����)�\��Y���:#���B-�q0��������eτoYF��R�(r�a��$u�	����:��j��� ���n��Cu�Eq��k仐.FN��hB�x�\O����[^Ơs�
\��m�RK�Y@E*�r�`솶������oAn���[g���r�@?�M�KZ{Ý
�OoJ:.�*�i=3�#W�2�)�x����KS��_:[(T�hV����ս���$��ӌ
[�ތ�t�s�2����4�}���:$^u��<��}�l�vk�P�����*�U�v�PJ2=e��(�<�$:�������)�俣��`h
�|n��Lo
m��[�h;X�ϰ+���A��T����!�cI�X�mk+ց$�|��@*��]SA��i�������B��� ��og�|�<���(a�&����w��ȳh4�5z����a�
���;R[��ّ} 5�N��Z�bV�r��t���%!�tf�I	
����Z��O����_>'��A���`� �Ȥ� ���Cfn����0�6�<�����[Ś!u�_{%p���&�<\%�K�����25�0�����GAe.��՘r4[/|In��=\��Z�b�����Sd��.��ﵽG�b�=�a�����t�����ob�S�qR�����F�=�p���?�HG���\M�|�߈e':� kBW�D(�ߦ���@	?��7��YF�&)�U��rA��;|�X�����|0�=�l�Q�~�т�������q��Jsk8��&¹���
V%2��(�%�����:��D���"k�&P�Y07������{���䟻�Sң��q>%��t��=�>��%O�v���O��^[A���?�d��r	�4ʉ���3I!��L� J�2��ҩ�Yh&R�(1�l绑���Ug����~��w�H.��Ov.���y�Ə��&EQDj�rCT�5�#LMe��
'�N��	�o��<V�n�"���mE���l>꺽T�li�M%����̥"�G� �s�5C�+E�E'j�#�����n2��늠Sn���s�7���׆
-DS�j|�S��0��m� /���E��= �}Q��.�.H�mȚ��(r�]����L�^r6P�弳��NF�54���K;��W���cV�g3�����m�y׉��ޙ���pj{�"#�i��/GD�a|mwj����;�oX�m�h;�Z1^�B���|b�d��
�������&uD� 0e�)X���~�m\T��rl���B���ӧ��u�d]p����z������g�8ӹ���]�Zwh$q� y�INa� .?17�i���Ҷ4ĕ�C�}�/����ޛ��n��<�V�>��^�:��=��C�J�qsN�T����fK���瞺�Ut">�M�}]��{6u\U�w:��\&�ڹA~c��$|�S��^F�4�[=6LN=�bpv��~b·��O�hd��&j~��w��e"�}kQ#2;��t��]��?R��2�i�A���+��`�j���Q�u�e�r�:b>�.�thu�B��|�`�Xq�(ʾ�n�f��H��DA�G�QV�MU"�8�bH��\m֡٩k�n>I�>IRx�{�d����Tx��
�#ԎLa)��'|���L����g?�ֈ����_�A�l��=��5u��X�4��y�4��i��s�#Qz�� ����qBBUE�]�ԽͅjM�g�_2!A�"���o�SY-��V3w<c���혧�ͮ9��2��i���ܳ*��Y�;[U���ｄ<P*]|/�X �c&Po�/Zp��@XL
� p݉ܣ�l�S��� �I���cx.ELnU�vvf՘�[a����
���C�R�B�u�Q������������Ί�8�́�V��@�_�<����l���V�E���nʽ��s<�E�Nu�	?|;�T�l��H�%��J�YM��x�tE�Ё��R�N
�EZQ��OV����P���tw��G%,z���J8��e�^vyHp۞����x^��0x~hW"�`�ڇ|m�g��-}$�=�B(�pPb��z߻�C���5�Wl������,���c�H����F�����gW��$j��xg�r�HB
�����4W�ĝ2i<(�D'�ʬ���D�^�Er��ͼJ\t�z[�NY9��fm�G�7����������l5[��v��u�va�	ޤ�EL#��c F��=}}x*d�ԋ����#g��ĸ�s�?�� �s����J�� ������C!zK����*矼��_��r�8v�.�}��>�������#g&[��������m�^�Yr����P���2v͐�d��Y���C����"�3�e�νe+��Tm��.��g��~��h9����q=�D��<�x*�%�Tb�N�B��?G=��<F�A�g"o����}��o�wA��bҲ�2��8g� �|�HW�;��S��{�!U�ZuϮ��v\(�I�� |��>�����=K��_��Лi����uS]�zO�n�yy���u)$�*eB���ùH(o�����`�0��hE�9�Ow������v.�L��M,ԩq�9��KMw���S���~N���0��Q�b�9q	�=0"�t���	iZu�5�+!�������Sۙ"��_|Ov���#e�w�����'V����!�-�[8̓��*�Y�FmnQ�u���?����}چ��f���2��D��0ݠDҿ��mT�����9��>!�]3H]�~�4a��]Y\o��辒��>!�;A�8��j,���d�8�g�l˓��HR��H�U��*ұC�d��ڈ�Y#<��,d��߱<����Hښ*�S�f#M���{��L)��nѿ�G�ׄD�?���<�]��bo˨�A�6.�r��57�+�N�Y{ƫ�eu�	@�u��B�l��|Ԋ�5x��)�2�՛��\����㖌���v��Ʈ���U���5�"
Nb���<�G��4����r$4��[���s���t�U�;����w���gȠt����Э��G��C�镾fQ���Q*X��寙4	���~k�*�.曼�Z��@-)*%x>BWRI:E���3K�ߋ�*b A]������P�m�I����3Т�-�
�g���<B�a���HIF�p�3 ��q�3IIԣ'=��%K≯[b�tl̾w�� ���)N�A�RH��<c��n��.7:�?n9��$W�Y�<5�~[h<,�Pv��������n��Ͻ�x��>z�5O1n$_-w�R�
�ɲ>=�9ؖV�c;�6x�W�23��SϿV}�Q�������9^�[������6�*58��9ت6d�k���(��f�+�qі3/∬;U�c��N-�B���T��<E_��,}��fh��U���%TŲp��r֞w9tq�O��) e��|��
��j���{y������!��IY9;�O0�����vl;{���SCU�;�jl�hO�I리����+�~{�cFc����TZE�`]��XïR5pĎ�4�1��Y�����D���|��J�hU�d6�x7h��\�O��f�g0]�b���O1b��D��ݧ-�*q�r���[��?=�}�Z3 >Vo/;g����Rڹ�"Rá