XlxV64EB    1825     990��b�O�� ��z��EϷɪ��m�r@��p3�	7�aC�x#U���ջ�Rueq9Q�aשR��!
-$�H����)�T��_�F,�킀�61v�a�U��堬Fgg�-� :��쏮Gn�$
w�f�rz����mV�%!Wg���-�����P� ���D�R��H:�ڌ����K�����S�urƼ�sa#�4Q�]�`�oV�WV�5���ր*��rA��F�1KY%�
�1zPk��g�W]`�+m�Xf��]�7���D�ܭ�b|,�[~2:Y�#'�Ν*�w�A�n.�B�ɱ�	�AD>�4�F�e =����z�ґ񳭏��q��̤{4� 1�
r>S1v���<T��;��x������(sp��
����TM�u������ ���r�K�SS�w��fru2�0P���,����:�
�߷�3�=2a?"਀�nM�0%���{��id���DeqLӫf��V+��0ɱ��j>U�n�呩X[��$l�q�Ֆ���U3���Y��6S��J>�In^y2������H!_�ɖ��NoDp��N���7[�6aIK'_"��c���5�c�3�c�A��X���QH�jFsp�.}߶	jj٤�!�9��2�'j/�5�	��fwsY�'��Aw}��hȎ��M
�@�(�}�سسLv��1��?(��t_���H�c�G��w@P�Q��%��q������o鑽��W0V~������$�N�~H��0A>jHD薫���Q&��m�\:��#hϩt�1�h.ᐦr�pz���řvW�;#,nb�U6[Nw�6���u��G�&���}�T��ͤ��jj�S�מ_���1�l�)R�yo^�T�`ס �%�*�&�Q�p��j[	���ĉ��W��(�/��eZ��"�8��f�����ڻh�R�[M�T4%��
H^t�C��c�#GXi�l��o ��ga��D�%p�Q�f�k�z85~�`}�H�usw�8c�y��i���t{�<:�Rs�5&~� ]�#��=��g��/����Ѵdu���%��qfj�B��n�:xߕ�ؔ��(�8�iG	☂%�T�&:��A'!N��p�5*�3wiޏ��~/떢���k��^˹aA�o�
L�{J=�ʐ^��#�rg��|��K7�*��{p�4��|�3����QN��1�g8�	0��Y���@����P;Bx�V8�E��H�B��C`�K��� ��}4��x����eS�C�t'��Ƥazc����{��j�+��Q{r_�
���� K�p�ǫ��J�ͳ�cLd�8�[�~��|��w��N�M8te�̇��Ĥi	����}l�?z;$�:-�3����ǐ1�+9>x<���I�9Q���j�)��b��|4.(,�#T�m����E�Ch��C<���4�Y�kĖ���Ԋ�ؚM�6f�e�s���?Y�^EcIYo݋[*W` ���?kG��}r��E]�Z��-��ha�y )'3T'�6�c��o�5�-��?ۨ�]1��A{��b��#Y�4�tAl���p)b�I�rgU׳�%�W ���J�ېS�ݗ@��O9��k�봢ꭚ{oa�B�c�z�ՅTc�����[Y*ZHs�t���q�	h�Q(f-�<�.A�[�b�[5�	N\x˧ʯ��UQ5� /��=
- �����a�[�ĎѺ���U	;!䎔����t����<텶��l�&�HmԔm.�Z[�vZB��Tq��K�{�H r�u��ٙ����}6��� �j���Fx��م�������x�Ez���fFo��NnP�i~9����*p	n7��Kp2}�O�2���gVKqh(v�C?2Q>}��,t��U����}�ǂ[mj��G�L]�A�w��C� &+��r ���*������HM�΍@&�/Z:��U$gO�yȓ{ݴ� i|�1+P���[��.�㑤k#ݴ���+d������G���~�oO��R�.�������S�;M"�P���4!������5��z�R&���&��#���Qo1�ѐW��^�F�ۖ+�<ѭ:����ˣ���^
~���v�<����ɹI�:+���^x���^�}e+��Iq�:�t/�| �{=�L��<�R{dGUt�c�ˌ��p-:.�\�x�s4FuSEy�U$6��^9�1�ܟ܊�hLПdu�fC��[+��k������>��)�J�V%i���3�<�1v�1�j�",�sa6�@3��#kd��|�<)�,�57��T��aر6��ܪ"&����_���0��_�9�'f��E�~�[2�h�v��(+�6��Y��r�z�l|�v��᯸+o���ol�{�7Oԍ#j\2"�Qu0���]5v�]�qs]B� xq�j�l�{�P�w�