XlxV64EB    15d6     820��ј!*25ŷ���Y͜f£�SĹ&�o�v	;��� ���}my�~ۖ�x�n��[;�(�2�����Rz%������a?�ʹv'V�8�oiM�vZ�	�Y5j��k9��j�6 ��˭��%KH��w�ey����4ţ�jd�����Ŧ�AS����v��.C� j����m�}A9Q�N��6.*�/��N4�Ul�H'2����w6<���\�g���ƃ��$V�_9\�G�L�e{<�;�����L�N�Q��m�����}ct��)��/2�M�S�3��("������T9
yXP�K"�@"R�m�t d&3�����~m����H"�^�N����Ӻ�y���/�a*F���]�{;jE0P�G*M�\0�//m��*�|�҈�qM7�V�^�f�5Д�U�]�T3��[��E1��>IΣ��K�v��c=���/#b�Cw��m�۟u�u{cLgBz�5�ʹV>��}�����w��i1������Җp�&$w�a�3WPo'��X���iQǘ��Z�F��J�Z?�	fTQ���0׀[ �Cزs�Z:�Q��<l�c�[7r��w��D���`��ÀgS�a��ŧ,�����qZ�֕Úƅ��Ix<�	�Yg4X�3�br��c,�3ŗ
�z��p����6�B_�Mf�*I��~��u_�#$�Q�L��8���wA�CJ B����q+�e�]��h:T`[>f�Y'�wy�6͊��q4ɜ�U���E`��ߍš�	Tm����̓����W{�����@Vz��_C2�w�&޵l��T�Y;%>ɹ��F4��A�����y�<V��O�T�I���� bӆN�ɧ Ei�c�@���!�!a�QKu{���Ɯ��*�Ox���o��`���JH�-�%�[�0ߋ���6�Dve`���N���Ħ �5�1.i�G	�V�.=2>��M�|7*�t�?l��J�e�g\o�'̱���3�����ǲ�Q����%�(��u�>bz�=^U���.r� �1U�c�9u���3V�X����;�z[�}�� J.�	�)U��l4���q�6���S��j�Lq�e�33��շ,�caaª��mL<����ɔO7�7�p�A.������t�=jJi�P�'6!����q�W�GZ����֡!:�);8G,��<��}.Ȃ�@	�x�Go�Rt����ka]��eJ;��cq���6���=�h-�e`���1_��G��[ʔ�gŞe���OG�$g�[�������G˱� ����Q6�P_x��d�w�^�?�	it�l��N~8Պ�y�A6=<7�5�Ɖ��G�wY[Hx����gq�f�Vu�sc�y�,:!ͽI�U=�.���o�}���s�lEÌ��G��a�ڕ��v�ʻ�q���R�6�&��J�I���PY:)����"[:���M�Y��Z���XM���X�ܻ�8�h�Jq)>6���O�Z����_po�<�ʒ�$z��e���6�e))��K�˿Y�5z(�F�4�
�I���V���e4ΉUI|#uq@�
AG���� >1�Qq�_\�GV�A�~�����|���nxMh!dbo�'<V�����F�0J"�5f�������������,Aj�R�巢���BQ�c�S��7N���CP�P�ߥL�xa9���P���γZ���C�p����2��K (�1�̫����^hG�l��L���z�/*������}�PE��pA���E�eFb��9 �o�ko��?|�3g6�+_5N�~�8- /��[K��G���r���Ļ'����h'T����$Z�g�^��y �'(��l��Q�s���$s�6�A��DL����p��({��ǭ�kB:r�ݬ��־e=Z�S!cJD{��M�QFw��n���Zo�7�B�k�Dy����e݄��b4ta��!��κ
�Ѭ��I�ң�.lV�YiZxe����K��C��U]����:A���֗�[�(n@Ǆ;��P�Ä�`��*�
��7^���x