XlxV64EB    1928     9b0����n
ղ�Z���a�t��Q ���#�P%�!>��������.����R��i����7ıcblz�z�djjz��U!w�1�߄��p�9��o�m��I���6۪ȳ���3]��"�t&Ŧx7�I�Ѣ0��)�1��k��)��g���%�Ϻ~�
��������N)1a)u���N�b��(w1�D������u)V�����5���e@���]�6)����&��(=	1���<�CK�A5UM��9�/c\_�4� ��A
������w|�;�3���c�`��}�-��]_�O�t�J��ӧR1��R~�V��]���4��
L�n�#�[�����D&��B;L���'�������Jaۜ��"m����3d���֓o^�4�j<�_��.i��M'(>2Ny٘�ϠL
VA�ҩ��i� ��1I����8-$2���� _T'�wR��i_�S%�X��'�;�SO��g`l�S�N�.����圄ձ��y���m�]g��<p(�RAOC��(�8hXo�2,jw�Vt�F�]�i�{s	V� Uoy�B���[���3�1"�r�U,��1�j#�E,wB�[s�f� F��A�q�K�_S/7V(ㆩ�}v|;ɉ�-�O�Q��;F�RBgE����|����;A��K,cC�P��j�k]
�ݒ���,F�a�2U�<�;O{�"9�����:_��+�!{��)ct>t��#�V���e]�h�K�m}8�����9��?�����&cU�ٸl0�{�1%�z��"2��[��O��zO,_%v뱣P��Y���/��ɩ����H�a�9�����KT���u)�� n�_�p��������k´SG�~`d��y"(�m-���1�'�x�9�)'���nm��j\{�u��`��U�.X��B��BI�u�xd�`0�P�>g���}?�#AQA�X�d�f�����0��1�L�P\)o!��#�P�x��٩P�����nʂ7w�Bz�*��R�h|]nY�����f"�Q�Mgz�r�����jK�W�εw�ɳ�,�	��"U����f�
H縌(��Лq���h^c���e�Gu���n4X}ά����6F�
ި�h��C��_;f�y�
$WDI �B�'�O-����8_}C� �j3l�t�<m���K�0���-�����5ozg:���@���
j��� �sS��o�V�o{x�Pgh\`�3.��`K<$mK�z9]��Ժ�Ŏ�?�:U�]�K\���Eu���b�@A�Ȭ��/`ń]2<���? |tȣp�����g�y!/|>_�*�F1��sJT�[�R�n�AWM�tuv��@�Ӻ9D�rP�}g�}d��$��ߨ�7|ˠ�ݨne�C��Q��bW�C!|�Jn��#�^n��bz���w���ع5y�Პ���y���B���g;Z>��WDܐnQ�O�t�̪u��ٖZ|r\ӝ&��&/t�9MX�0O���EF߱�E�^��6�V�K�^��0�Za	��J��{��QG~R��I��D�2���0�LO�	���I0�J�y�dB�߾���l���j�#����:�sݻf?�Yr}�{��>�ģPV��o�j�JZd�.���=�t��߰�����#�|�V����b�iz̵����@)ڜ]qC"�pY9x��ү� �fa-�j3蟋{z,�n�����	R�FO�Xgԉ�!�1���ey��V�M����R��}v�v+W�x6q���l����=B@�ށH;7�-&ĥM���pbd'?ݢk�m����x���9������<q��.�!��O�pg�n�\�v����K&}0):���&��a�*<G���x86N,���$R�o�٣��7�5�%��	2	�i�TJ?5��u�-�z*��⮝l����r
ˇ&���η����N�¤������Knƀ1a�M��ȯ�Cb���#r�G�fF�%'�R��Ġ�*��y����ZF�B�5n|_9��Ӧ�[�ti,AB�n^�y��W Y���e�Ǜ�ʟ�U�c�X|�r����ȿ�@^`|@f�GD
�����2��F
�ê�reգ��d�$��uO���)�1�	TnM�]�s�]J�׼V��Bi�HT��4����q+�R�O_����U�Gl�o%Ű��7+װ�w����a�����Pg�H�_ڪ���A���i 0��u啳�#UK��'���l/���<�O�5D�P�s�"��F�c�>�m�`

���حY﹖U�|�X�9d��~�V���B�_��I�!��W�~� oe��z�����Z�՝_��(3-3�܍�<�_S;���0�u��.�=�Y��8�PO��-]��������V��ћ����v�$��!�T��(m���^����܎��M��d>w��a��|~1