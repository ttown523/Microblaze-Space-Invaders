XlxV64EB    5743    14b0L�/��v�F6�PRQ��'eyK�׉̭gMeΥ���$Z����� ��?,?�?���!��}��߿1��j�ýݛ"(\����?䔛2ItHɱ�#�(�ESO�$	��^n�m=���n�������O}k��
��B������)7'(N{M��aHE��%�j�r�g���k��{z���${6�l�U��$��O�������A r8��K�̯�@���C��]�V�����l�v�O(�8��	H	�5�\ԗ��첺����04dnz���	�+�.�T�}�%_F]a��x[���u�������U��_�����Y]k�<��d��;D��
>�#�pm*�X��#g��9�1#*9��2cw�훌��!�6y&z�@Xg��B��Q���?��sy"�6
���0��Cg�Nb�Fk���)IP�8���^����p� #y'Cԡ��#pcy6r<��Ux�,zld����4?ݫ���oA1X�ݱ�TsE/��[R,$R�8���BWj�Ȩ�?![dK��$BڭI��Cy��e̟b@>G���4���l:��0�:�.O��ْ�])�y�n-Eք��"��*�ю�����K�*��}C��������=%RB�:��s�އ�����
Xl��I:3�3�٥�*(�D\/M��Z�h��JV��^-	���;.��0Gq�R�R<U
j� I^L_r�JCO��>X�r̗j��$�pĜ���*�5�t�v`Ź���X>�$���~��o_벚A��R��(�f�=l<�V�����x�`����,�,�c�_�S[T���o������v�~��P�'r�/�iB|8EDj�o9������}���e�y��#�V���XAD���]���ET���u���������]$ɕ�%�"KK������*�|����-�t�|��)�7��4�?f �)��6��ٺJ�u�g�.����H�+9n��V����z��L58�6�k��M&ݲ�Mŕz��� �N{�Q-Si�����-(iF6)��b��8��с.�L�O�
o��5	�:�!8�.r��aQ�����z�k�����C�ثG�g�׷�A��Fo��'��p��q����p�����2���߈�g	�g��+ah��ec����ki5}b��y�}��|��f"ylI�M0�y6g�ݒ��]�ZcJ���I��>q���k=t:	{�^���&���<3%YgTv^مg�7�^��B�e&���NF~��ܨФ=Ŭ�eR�t6c:�Z7gO�j��mQnM"Nv"G��N�[8�u���w���}-�ۺ��ܺ�b����@9���?���fiu*��>٢�1�l�����^ߝ�y���E-�Gdh(�8�gv�.:[턪)N�o}��!�2C��:i�m�aOK��������3�a�9s��a��Q��ޠ��)S�3�t� ֮2Kb���Isl�N�̋����
�'�Aw|�����(;�t�Q����D�0P�	w�������:�I��Ԋs{�6GZ�(���D4{/�g�s�e&���crR��ǫoU���Z�O�4�-W���L��u��(AY�P�u9�2?n'N#��hcs��JsE]��5z�/��>����{���KZ"�b��#���^R�ߋPdŶ�Ťc>ұ'������@S�S�g@��@��r�=躐'�IQ��Ei��<~��� �>(o�}G� 9�e+qPZS��V{_dY���4 ���!��_�ޚJo�W=F��ɅU��
<y�&:���Ǽ�r7Ζ��ڳ�J�ͤ��%�j)|����DZ��N���,��|6�sy E�턐o!���^S�{��ʳ�����2U�li���WV�z�dek�M�����d*pNR�����6Cdv��#(��u�!fo���4��FN���#���ф�]ۂ�R��{Eb��+Г�I�����湇���������s����ȁ �����y�oJ���ήfk�+/��-�/潵��d�����&I�$}��-� 5��Û��_s���L�M��4x쳹J#g�s8DUWkL��p��\�f�jF���A�-��ΔD�����tZ�}<��3����Hb�'^䝕�^�(S_ʊ�퍭�0��{2@��������-�|m���a�?��B#�o�sh*?��.#f�/&�I� ��VE3�T���L{��m4t\��]y�E�V؊r)��#LR|c(�w��[��@���|�ئ�����y�OU,��è�����jmQ�3�96�ksH��7y_��ɡ��D�ݕ��
��e+D��qGc�/i(��E��*�$�U���tvH
I&��Ԋ�T�b��#��w%�h�!���[��ޟނ�..?��{�6rՕ2c���0�,��!%P���E����(����F�s��T���6hdz�c3��$�[�)�FrD�${�JUm�4�;�j��� 0P�m�b&J�.K$_ qh�E 	�s�1h0���d���y����WB��X��r��W)���myج�'�hw��Iī��E���}zI.%�4:�0�I����t�6u3��˾!��^F2z�-@�.�`��� S�S��GV	E�z���@YE?_��<y\����<D�����2�r�o	�kGP1cߊc��b��P<ŝ�Y�Xn�Z�����X���]un3W�B\�A��Ŝ�-�U[��"���.Z�
�V� sf�=X�ww��v��%�
�~3�gZ�t�Ę`'����O�(��G����dHq�p:/#�"_S��d����ʴt����՜����;hlK$����㳚�'�U���~�͖�,UKyı�z�5��n�ą!�g59�eFŭ������K����D�V�O��H$�8��q�ػ�A���5�8�k0�����_�m��T�}t�<����r�8;�A�G�D�Eʇx�D.y�#�@_ڇO���/��jxY��o��g��c�п�_��G,�;�(4D��_�œ���^=��Or4ӛ�#�IΣ�2���*����:=�C�QB/+�$�k�n�����]��W�۰�I�y��uLA�n���������9�ҳU�PWjp��3����:�f�Q���+�]��EgV����#�X�:�����qŁ��-��X�W~�^��y'ɟ�k��W�))s�-���.Y�C$���?(��� hѢ@	��Y�3W"g�j �{x*����d�ƍ��5�0f�D�@�'#a��5�,��H9�pl�W͒�1^�������Œ�,�v5�p>]�#�*�������^�s�k�R�Ѵe��B=+u�����`�ߧ��&\�����S��e���t��D*ZN�#�d �O�#J�喓�a�M/>��:�g��l��V��a�!���k����I}�҂�'d����(b�@��Gb�'��h=)������2x �����c,B��T����g�V��b�8?R�sr/L�ݬ���l��F[�� :��P1���Dʃ lb'{A�����*��*�e-��$�+�v���޾gMe[�,��"L.��0]*D�{�&�������*Q��k���[;��Y��@��8�J��qX�����N�P�%��J6}S�}���M���͐��a��xL�9�B���sW^Eo�L����1���Dq� e��A䲇�C�����?C�3-*��)��0
}/����_�XK�؏���0��M���%�^7��cg�4�C��&����{�\�ḟГyFQE�Y���e�ՠ3^�	�\t�b(�Ywcofv ������KT���Yr��4��Ys}�R��h	�a��H<��:r�P��R3<����Mx-Hl}A�0��yap� �H��y�t/l����޽�e�3!�Ґ>n�n�I��r]��[���n3p{�O��SV,uv��>�1�9������ߧ��o���'[}��[Ua�?��1`��x&z�ê�m!ag2��B�{�6�n-���d#=)e$��"5v��u쯠yh��=?���'��\A�e=*�����^�h�K�ڡk؟>.�#��z+����*a��D�$#S,�i8:�g��|���.H�J��G���4K�oj��N�o�����$�OI
&((& �=��y�e<�o02q@�`N��3}��|DR/��Q���U�I�a��Y!z�jD!�B�F2�H�*�D{�SS�;6}⛒��;�g,�ɛÅSL��	�cF������T!B������m����pє�d[�]�e���C�� GBY����DsT;�هAD�-'֚�ФXz��S;�(I8�P2��WbO�֡�[y*��l��K��$�nC:kx��]�����mF��������--�Xd�Jj�l0�g���`9Urm����K�\��l����[�Q:)Wm��#�]�-��-���_�X�+H�M����F�F�*��)�RV�i]s�v%n6r���k:.6��ɂ�gJ�L�A������+p�q�hm @�$Oi:��B>q,��$�>R_��z�t��i������f��%��'�����k��#���ld}��spM��h����+��܆4Ӳ<��]�K�jL����}V$��rH���
��Z?�z�������?5�4N��cU�n%�Y�h/N�穀��rf,H���u��3� 5Ղ�lr%f���~;�`b�F|Y{�~sr��LIOmș˿@���~Io�ic�E�a�J�֐3���)сz:� �s���<�R��rP샓��"�����1�����5�C��ͥ�g����a%�)M���[���r�"T�~B}h����ro�J��[}�b�%TF[C���R��8\�*�`�z�CIj�ğ��?,r��*� ����#����L�92�%9�&�&�m� ���#[�����X�@���¢�f�� ���ݙ��!|PHqbQ�~̵?�\$�˜�-��!�M||�6h���e�G#5��7��O������!��H�R˒�(+�B f�����BZC��H	m��Ѿ`�?t�-���-���n��/~�����R��Cy�<���h�ײ�93�r��h-�.���Yf)��;���E��%�t�
�u�Q�
�8{�_���>���g� +:�z����o�!?�xXxU��TR������F��e C�N�9��X��9���:\=3;��(�J.!8#�*^��6xI��~�