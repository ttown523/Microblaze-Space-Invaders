XlxV64EB    1554     7f0����S�A�E�&0{�W�5R���B��Ť�v?G	�fW�f=�+7��/N%2ܑA*���%�Uz�+�һWD]�Jb�5b��T��1�W��`�y��ë��!F���kx�ι���!U��]U��)a=Me�'�XMo�Uz�o��3x�7Wg¢4Q�Wo&�o��8�]	zi�N�J����\�]��_�T8��w�L��̯�obn"R��΋�Q@%k�ڴ+~�g�3�/��dl؇f0���Zۃ�e���C>?��4�u�j�q��w�𓰪��{����IB9'87d)�N5�4�;{%��?���R�Eb�u�+hP��Jyn��z��G�ܼe��:h�����_L���f(R�wV�H`�w�X�4{&�4ё �V�� �2���,�蒻�K?˖)iϧX4�B�L��ݟ�\x�5!.�kȬ��LW9=k��(����P|����EǊGu"���Gz�I`8v�����p��hi/A\8J�F�r�mB�d�C�Y����(-�U��	�a+e{��-'y�}��U؄MI�(�˫E7�28o�xEs�l�9�,$�g6̥zO��~�9T��؎M�:��s��ޖ
ۜ�?7h��c�|�Q�kۺ��[����t�n?C�,)�j3*�O� �S��;fd�b���}\��GH��v���g�]c�vm�����Y+~xP��]���?)�zO��n6��K�;�V�q�\Q@���Q4|�C��*���3�¹u��}lno�U��.8�68�fмȰ�>Q2Ї"`F�����/)�t~pʏ��,�Wʥ�IOUXu����Y��Ss�k�1꺋T��mc�r���	Ό��v5���f���?�-�}����ȿQ9X�K���>�k�� ���iJ{)+��r(��t<!�����6��w������S��X��3�d/]q��Gg&���4\��߈�p�8k�Q�,f��1��o%���������9w|iy҉p�mf� ��}��̜
���1��G?q��v�8г�:)�I�^ɔ}Z�3�n���Ӝ%��	adc�������)�?-��5�{�Y�%���#>�?����*���
�x2Q[�)��_pm���^B��ٞƽ'�����)�K�N��֒��A����=FEA�֦�<ӈ�`�
ٳ��E*r��٘�Ů�+�����rQ�Q�g=5݀�`H#q mч���Z��x�r�sYK.:66�����YYX��+���V�+���Q���h _E��܏9�~���m��a)J��tP<xO��5?F�?���0_<�v��<$��<��fsǙ�`�4z��4B�����O$ϩO���?�2��!����X�
I�u_I�&�����(�rGXݥ�+l��ٕX`���
�*�B*��:qؼK�A�ǋ-v�,�C{�{�׌�����N�4��(IM�UY��6)�i��X���CЕ��~n� �Z�!¨п䦸����\Ga�B�i����}Z`��S�K%�WEGJ��
�r/f�����w�`P���Z����R�V��(�~}7B�V!Y�
���.
(?dl gn��(1�l��y��U2�����0pܬ0%FJ&��?��E�� v���*;���2��#4��N�+ޢ�@>�n[V�'����ٽ�u�w⏛����i w؞�
���􍊦��Gsv���p�|'S�U$�3Q�I��ԶW�A�aw�T
f�&B$�A�Wy�@JA�%H� ��t�$�$d�x^� L�'U�L�����F������Z59�$�մ	��?X�<�ܾ�|�R��6�,��%`^����(�neN*z��N$�)4�п�'���ZZ������I }{�߻�7�v~�A���d�!�7�w���H���.��)3�_�X�(�T�մcA0��r�n���J>��F�'�&;Ź��R1�����5p/�茞��vvZ����"�V{�kPn||P�¡�3[�?�3�[g�{	n$����