XlxV64EB    1846     8805��8R.:���Hkȥ;7���Q\И����ȿ`^��]T<��.<����,��d]�^}�v^�w��_��4�i?��A+"�:ʰ_�;�'U�z��&�D>�</�z�{�,9Xi"��P�UIgY��z-H�����D$Rbʌ)�=�.�5�	��h�W��&zg�]�f�&�A�8X��˰�}x�E�t?����~�V`�D"!Ůj.���!����j8������I��pg$�*۶u����:��47s& K)'��G4pL��g�εmx�Z�`�8��@�c��z�L��劊S�Q�t���!�F�M=�>��m��^8o���}(⾊,�_�Z�pC�lB_ΤIq�9g��.���h�K[���P3��n������δ�[��+����͍ V��By�䋃.v�N��C���������	$z��y#U>l�x��+�N�&_�l�S� ,>m�)��A�ƶ�~
�˔�m�Ϝ$s-q&ݳ0�,��Rt�]BzC�&6;M8��ɕx�����[�ʡ�l�]5'Ql���p�37t�D�ն1v0a�w���U͓DI<�WTc$�#Ny�e�ƽ����H�n5�`�D��B?�s�3F�^t�{v��o�-I��B��1k�1H ������)OפZ2Źx�%N�r����h������}�~ |+hk1�&!�rQw Pf��y�O>[1�h �>�g%Ҙ65�����o��3���j���������Ql���ot���#^�P";�g[�2LVYm`!|XK����H����}`9����M6�;m����ݛ'9�C�(J�
:3�e������x�>��m�/�˒(E˕�]}�*!��YI4��� �����z �k8fr�+H���F�N�S�L4���N�9�4&M�{|J���>#��"m�����I�y�`9��0ÁL�?�����&����!�4d�876b�k�u�K����s�؞p��4���ʒ�����B�i��Y�s�+��ޙP�<q��볗��=>S�o�d�I�ߞ>شGV#��znJ
�7�F|'����$F�2�%�Kx3�(S虄�ٳ)�WCP|><�b=��A(�]�q��z�?���j��SG�bl-~���&�lUG)��՜��C��@"LVP-KS`�[��i�0�����sg�v���L��:t����/.&��/�S=F[�)�G��*�:v��a��m�������sF\W����o����M6;Yu���4c��B�Ɗ�7��J�����p?����=�B��
�aE�J�e�q�m�{���m����n܁pZ/�J�-m߼�G={+>�{�oݼ���ܦ�;�k��w���׋���ؑ}�XS��X��_�h��g��y���[��{�
���(�4���6�w�2Ҩ;���;����⤲_E���]\\��lu'�6x�#<2��]�l�����a�R�;mX��fP�aX$n��I���cr^��=Ġ�F��( R�79Ժ7]�:(��
P� ����k���iOğW�6�$&��dZh,;<3Y��
����6?��
x�,��81~WQe6��[�&�g ��:=��F�8�s4���E���1�s���3�z��K��LU���APU��V�|҆GV��;,\�_H�N��QDt�_Ciw��=w���M�
��C��6~v9�yڱ��)�1
��%;�B�z�dx�	���`W0�g��"���Sf�ҭ���T5��}T�(�գ��.���<�W�����}ނ�F%%~*he���O�g򦐍�E�5�Ec*���4��CF���F��"ټ4!��пLs��a��,���Iu� jͪNY��U��������V�_�ڀ�jO�&�KS�|���b}��b,�p@�2$W߇?���/��PK	�]y(	�LS��)�R��/#e��a��o\B�1����~a٬������CC\C+���m�����tw���w�	�5���$f���#;1rcs- �/��P֡=УQ���ߺ߳�X�X�okhY��*�	�S� �����\v�-R�������ʇ�!��P�T���4�Q�M��_�^iU��}+`����ݤnL��,���:�����@���D�N�|?0���|�